
module CTRL ( clk, rstnSys, startSys, rstnPsum, rstnPipe, rstnAddr, addrInc, 
        latCnt, start_check );
  output [15:0] rstnPsum;
  output [3:0] latCnt;
  input clk, rstnSys, startSys;
  output rstnPipe, rstnAddr, addrInc, start_check;
  wire   N17, N18, N88, N90, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n3, n4, n5, n6, n7, n8, n9, n12,
         n28, n29, n30;
  wire   [1:0] currentState;

  SDFFSSRX1_RVT latCnt_reg_3_ ( .RSTB(n38), .SETB(1'b1), .D(rstnSys), .SI(1'b0), .SE(n36), .CLK(clk), .Q(latCnt[3]), .QN(n12) );
  AO22X1_RVT U17 ( .A1(rstnPsum[0]), .A2(n16), .A3(n17), .A4(n30), .Y(n43) );
  AO22X1_RVT U18 ( .A1(n18), .A2(n30), .A3(rstnPsum[1]), .A4(n16), .Y(n44) );
  AO21X1_RVT U19 ( .A1(rstnPsum[2]), .A2(n16), .A3(n19), .Y(n45) );
  AO21X1_RVT U20 ( .A1(rstnPsum[3]), .A2(n16), .A3(n20), .Y(n46) );
  AO22X1_RVT U21 ( .A1(n18), .A2(n30), .A3(rstnPsum[4]), .A4(n16), .Y(n47) );
  AO21X1_RVT U22 ( .A1(rstnPsum[5]), .A2(n16), .A3(n19), .Y(n48) );
  AO21X1_RVT U23 ( .A1(rstnPsum[6]), .A2(n16), .A3(n20), .Y(n49) );
  AO21X1_RVT U24 ( .A1(rstnPsum[7]), .A2(n16), .A3(n21), .Y(n50) );
  AO21X1_RVT U25 ( .A1(rstnPsum[8]), .A2(n16), .A3(n19), .Y(n51) );
  AND2X1_RVT U26 ( .A1(n22), .A2(n30), .Y(n19) );
  AO21X1_RVT U27 ( .A1(rstnPsum[9]), .A2(n16), .A3(n20), .Y(n52) );
  AO21X1_RVT U28 ( .A1(rstnPsum[10]), .A2(n16), .A3(n21), .Y(n53) );
  AO22X1_RVT U29 ( .A1(n23), .A2(n30), .A3(rstnPsum[11]), .A4(n16), .Y(n54) );
  AO21X1_RVT U30 ( .A1(rstnPsum[12]), .A2(n16), .A3(n20), .Y(n55) );
  OA21X1_RVT U31 ( .A1(n22), .A2(n24), .A3(n30), .Y(n20) );
  AND3X1_RVT U32 ( .A1(n25), .A2(n15), .A3(n26), .Y(n24) );
  AO21X1_RVT U33 ( .A1(rstnPsum[13]), .A2(n16), .A3(n21), .Y(n56) );
  AND2X1_RVT U34 ( .A1(n27), .A2(n30), .Y(n21) );
  AO22X1_RVT U35 ( .A1(n23), .A2(n30), .A3(rstnPsum[14]), .A4(n16), .Y(n57) );
  AO21X1_RVT U38 ( .A1(n26), .A2(n25), .A3(n22), .Y(n27) );
  AO21X1_RVT U43 ( .A1(n25), .A2(n31), .A3(n32), .Y(n17) );
  NAND2X0_RVT U44 ( .A1(n28), .A2(n33), .Y(n31) );
  AO22X1_RVT U45 ( .A1(rstnPsum[15]), .A2(n16), .A3(n34), .A4(n30), .Y(n58) );
  AO21X1_RVT U46 ( .A1(n25), .A2(n35), .A3(n32), .Y(n34) );
  AND2X1_RVT U47 ( .A1(rstnSys), .A2(n36), .Y(n32) );
  NOR2X0_RVT U49 ( .A1(rstnAddr), .A2(startSys), .Y(n37) );
  NAND2X0_RVT U50 ( .A1(n10), .A2(n11), .Y(rstnAddr) );
  AO22X1_RVT U52 ( .A1(n3), .A2(n39), .A3(n40), .A4(n26), .Y(N90) );
  AND2X1_RVT U54 ( .A1(n25), .A2(n29), .Y(n40) );
  AO21X1_RVT U55 ( .A1(n25), .A2(n14), .A3(N88), .Y(n39) );
  AND2X1_RVT U56 ( .A1(n25), .A2(n15), .Y(N88) );
  AO22X1_RVT U57 ( .A1(start_check), .A2(n25), .A3(addrInc), .A4(rstnSys), .Y(
        N18) );
  AND2X1_RVT U58 ( .A1(currentState[1]), .A2(n11), .Y(addrInc) );
  AO22X1_RVT U59 ( .A1(n25), .A2(n35), .A3(rstnSys), .A4(n42), .Y(N17) );
  AO21X1_RVT U60 ( .A1(startSys), .A2(n11), .A3(currentState[1]), .Y(n42) );
  AND2X1_RVT U62 ( .A1(rstnPipe), .A2(rstnSys), .Y(n25) );
  NAND2X0_RVT U63 ( .A1(currentState[0]), .A2(n10), .Y(n36) );
  DFFX1_RVT latCnt_reg_0_ ( .D(N88), .CLK(clk), .Q(latCnt[0]), .QN(n15) );
  DFFX1_RVT rstnPsum_reg_15_ ( .D(n58), .CLK(clk), .Q(rstnPsum[15]) );
  DFFX1_RVT rstnPsum_reg_0_ ( .D(n43), .CLK(clk), .Q(rstnPsum[0]) );
  DFFX1_RVT rstnPsum_reg_2_ ( .D(n45), .CLK(clk), .Q(rstnPsum[2]) );
  DFFX1_RVT rstnPsum_reg_5_ ( .D(n48), .CLK(clk), .Q(rstnPsum[5]) );
  DFFX1_RVT rstnPsum_reg_8_ ( .D(n51), .CLK(clk), .Q(rstnPsum[8]) );
  DFFX1_RVT rstnPsum_reg_3_ ( .D(n46), .CLK(clk), .Q(rstnPsum[3]) );
  DFFX1_RVT rstnPsum_reg_6_ ( .D(n49), .CLK(clk), .Q(rstnPsum[6]) );
  DFFX1_RVT rstnPsum_reg_9_ ( .D(n52), .CLK(clk), .Q(rstnPsum[9]) );
  DFFX1_RVT rstnPsum_reg_12_ ( .D(n55), .CLK(clk), .Q(rstnPsum[12]) );
  DFFX1_RVT rstnPsum_reg_7_ ( .D(n50), .CLK(clk), .Q(rstnPsum[7]) );
  DFFX1_RVT rstnPsum_reg_10_ ( .D(n53), .CLK(clk), .Q(rstnPsum[10]) );
  DFFX1_RVT rstnPsum_reg_13_ ( .D(n56), .CLK(clk), .Q(rstnPsum[13]) );
  DFFX1_RVT rstnPsum_reg_1_ ( .D(n44), .CLK(clk), .Q(rstnPsum[1]) );
  DFFX1_RVT rstnPsum_reg_4_ ( .D(n47), .CLK(clk), .Q(rstnPsum[4]) );
  DFFX1_RVT rstnPsum_reg_11_ ( .D(n54), .CLK(clk), .Q(rstnPsum[11]) );
  DFFX1_RVT rstnPsum_reg_14_ ( .D(n57), .CLK(clk), .Q(rstnPsum[14]) );
  DFFX1_RVT currentState_reg_0_ ( .D(N17), .CLK(clk), .Q(currentState[0]), 
        .QN(n11) );
  DFFX1_RVT latCnt_reg_2_ ( .D(N90), .CLK(clk), .Q(latCnt[2]), .QN(n13) );
  DFFX1_RVT currentState_reg_1_ ( .D(N18), .CLK(clk), .Q(currentState[1]), 
        .QN(n10) );
  DFFX1_RVT latCnt_reg_1_ ( .D(n9), .CLK(clk), .Q(latCnt[1]), .QN(n14) );
  NAND2X0_RVT U5 ( .A1(rstnSys), .A2(n41), .Y(n7) );
  NAND3X0_RVT U6 ( .A1(n3), .A2(n4), .A3(n29), .Y(n33) );
  NAND4X0_RVT U7 ( .A1(n28), .A2(n3), .A3(n4), .A4(n15), .Y(n35) );
  INVX1_RVT U8 ( .A(n13), .Y(n3) );
  INVX1_RVT U9 ( .A(n14), .Y(n4) );
  INVX1_RVT U10 ( .A(n36), .Y(rstnPipe) );
  INVX1_RVT U11 ( .A(n35), .Y(start_check) );
  INVX1_RVT U12 ( .A(n16), .Y(n30) );
  OR2X1_RVT U13 ( .A1(n17), .A2(n5), .Y(n18) );
  AND4X1_RVT U14 ( .A1(n25), .A2(n15), .A3(n14), .A4(n13), .Y(n5) );
  OA21X1_RVT U15 ( .A1(addrInc), .A2(n37), .A3(rstnSys), .Y(n16) );
  AND2X1_RVT U16 ( .A1(n4), .A2(n13), .Y(n26) );
  OR2X1_RVT U36 ( .A1(n18), .A2(n6), .Y(n22) );
  AND3X1_RVT U37 ( .A1(n14), .A2(n13), .A3(n25), .Y(n6) );
  NOR2X0_RVT U39 ( .A1(n7), .A2(n36), .Y(n9) );
  OR2X1_RVT U40 ( .A1(n27), .A2(n8), .Y(n23) );
  AND3X1_RVT U41 ( .A1(n15), .A2(n14), .A3(n25), .Y(n8) );
  INVX1_RVT U42 ( .A(n12), .Y(n28) );
  XNOR2X1_RVT U48 ( .A1(n28), .A2(n33), .Y(n38) );
  INVX1_RVT U51 ( .A(n15), .Y(n29) );
  XOR2X1_RVT U53 ( .A1(n4), .A2(n29), .Y(n41) );
endmodule


module OSPE_0_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_30__0_, ab_29__1_, ab_29__0_, ab_28__2_, ab_28__1_, ab_28__0_,
         ab_27__4_, ab_27__3_, ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_,
         ab_26__4_, ab_26__3_, ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_,
         ab_25__5_, ab_25__4_, ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_,
         ab_24__7_, ab_24__6_, ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_,
         ab_24__1_, ab_24__0_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_,
         ab_23__3_, ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_,
         ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_,
         ab_22__1_, ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_,
         ab_21__6_, ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_,
         ab_21__0_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_,
         ab_18__9_, ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_,
         ab_18__3_, ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_,
         ab_17__12_, ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_,
         ab_17__6_, ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_,
         ab_17__0_, ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__23_, ab_1__22_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__31_, ab_0__30_, ab_0__28_, ab_0__27_, ab_0__25_, ab_0__24_,
         ab_0__23_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__25_, CARRYB_5__24_, CARRYB_5__23_,
         CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_, CARRYB_5__19_,
         CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_, CARRYB_5__15_,
         CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_, CARRYB_5__11_,
         CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__26_, CARRYB_4__25_, CARRYB_4__24_,
         CARRYB_4__23_, CARRYB_4__22_, CARRYB_4__21_, CARRYB_4__20_,
         CARRYB_4__19_, CARRYB_4__18_, CARRYB_4__17_, CARRYB_4__16_,
         CARRYB_4__15_, CARRYB_4__14_, CARRYB_4__13_, CARRYB_4__12_,
         CARRYB_4__11_, CARRYB_4__10_, CARRYB_4__9_, CARRYB_4__8_,
         CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__27_,
         CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_, CARRYB_3__23_,
         CARRYB_3__22_, CARRYB_3__20_, CARRYB_3__19_, CARRYB_3__18_,
         CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_, CARRYB_3__14_,
         CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_, CARRYB_3__10_,
         CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__28_, CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_,
         CARRYB_2__24_, CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_,
         CARRYB_2__20_, CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_,
         CARRYB_2__16_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__0_, CARRYB_28__1_, CARRYB_28__0_, CARRYB_27__2_,
         CARRYB_27__1_, CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_,
         CARRYB_26__2_, CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_,
         CARRYB_25__4_, CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_,
         CARRYB_25__0_, CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_,
         CARRYB_24__3_, CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_,
         CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_,
         CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_,
         CARRYB_22__8_, CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_,
         CARRYB_22__4_, CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_,
         CARRYB_22__0_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_,
         CARRYB_19__9_, CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_,
         CARRYB_19__5_, CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_,
         CARRYB_19__1_, CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_,
         CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_,
         CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_,
         CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_,
         CARRYB_17__12_, CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_,
         CARRYB_17__8_, CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_,
         CARRYB_17__4_, CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_,
         CARRYB_17__0_, CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_,
         CARRYB_16__11_, CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_,
         CARRYB_16__7_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         SUMB_29__1_, SUMB_28__2_, SUMB_28__1_, SUMB_27__2_, SUMB_27__1_,
         SUMB_26__5_, SUMB_26__4_, SUMB_26__3_, SUMB_26__2_, SUMB_26__1_,
         SUMB_25__6_, SUMB_25__5_, SUMB_25__4_, SUMB_25__3_, SUMB_25__2_,
         SUMB_25__1_, SUMB_24__7_, SUMB_24__6_, SUMB_24__5_, SUMB_24__4_,
         SUMB_24__3_, SUMB_24__2_, SUMB_24__1_, SUMB_23__8_, SUMB_23__7_,
         SUMB_23__6_, SUMB_23__5_, SUMB_23__4_, SUMB_23__3_, SUMB_23__2_,
         SUMB_23__1_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_, SUMB_22__6_,
         SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_, SUMB_22__1_,
         SUMB_21__10_, SUMB_21__9_, SUMB_21__8_, SUMB_21__7_, SUMB_21__6_,
         SUMB_21__5_, SUMB_21__4_, SUMB_21__3_, SUMB_21__2_, SUMB_21__1_,
         SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_,
         SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_,
         SUMB_20__1_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_,
         SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_,
         SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__13_, SUMB_18__12_,
         SUMB_18__11_, SUMB_18__10_, SUMB_18__9_, SUMB_18__8_, SUMB_18__7_,
         SUMB_18__6_, SUMB_18__5_, SUMB_18__4_, SUMB_18__3_, SUMB_18__2_,
         SUMB_18__1_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_, SUMB_17__11_,
         SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_, SUMB_17__6_,
         SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_, SUMB_17__1_,
         SUMB_16__15_, SUMB_16__14_, SUMB_16__13_, SUMB_16__12_, SUMB_16__11_,
         SUMB_16__10_, SUMB_16__9_, SUMB_16__8_, SUMB_16__7_, SUMB_16__6_,
         SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513;

  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(SUMB_27__1_), .CI(CARRYB_27__0_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(SUMB_27__2_), .CI(CARRYB_27__1_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(SUMB_9__3_), .CI(CARRYB_9__2_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(n199), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(SUMB_7__4_), .CI(CARRYB_7__3_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(SUMB_6__13_), .CI(CARRYB_6__12_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(SUMB_5__12_), .CI(CARRYB_5__11_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(SUMB_4__7_), .CI(CARRYB_4__6_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(SUMB_3__9_), .CI(CARRYB_3__8_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(SUMB_2__19_), .CI(CARRYB_2__18_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(SUMB_1__24_), .B(ab_2__23_), .CI(CARRYB_1__23_), 
        .CO(CARRYB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(CARRYB_1__24_), .B(ab_2__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(CARRYB_1__25_), .B(ab_2__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  XOR3X2_RVT S2_24_7 ( .A1(ab_24__7_), .A2(CARRYB_23__7_), .A3(SUMB_23__8_), 
        .Y(SUMB_24__7_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  XOR3X1_RVT S2_22_9 ( .A1(ab_22__9_), .A2(CARRYB_21__9_), .A3(SUMB_21__10_), 
        .Y(SUMB_22__9_) );
  XOR3X1_RVT S2_17_14 ( .A1(ab_17__14_), .A2(CARRYB_16__14_), .A3(SUMB_16__15_), .Y(SUMB_17__14_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_) );
  XOR3X1_RVT S2_13_18 ( .A1(ab_13__18_), .A2(CARRYB_12__18_), .A3(SUMB_12__19_), .Y(SUMB_13__18_) );
  XOR3X1_RVT S2_14_17 ( .A1(ab_14__17_), .A2(CARRYB_13__17_), .A3(SUMB_13__18_), .Y(SUMB_14__17_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  XOR3X1_RVT S2_2_29 ( .A1(ab_2__29_), .A2(CARRYB_1__29_), .A3(SUMB_1__30_), 
        .Y(SUMB_2__29_) );
  XOR3X1_RVT S2_20_11 ( .A1(ab_20__11_), .A2(CARRYB_19__11_), .A3(SUMB_19__12_), .Y(SUMB_20__11_) );
  XOR3X1_RVT S2_11_20 ( .A1(ab_11__20_), .A2(CARRYB_10__20_), .A3(SUMB_10__21_), .Y(SUMB_11__20_) );
  XOR3X1_RVT S2_3_28 ( .A1(ab_3__28_), .A2(CARRYB_2__28_), .A3(SUMB_2__29_), 
        .Y(SUMB_3__28_) );
  XOR3X1_RVT S2_4_27 ( .A1(ab_4__27_), .A2(CARRYB_3__27_), .A3(SUMB_3__28_), 
        .Y(SUMB_4__27_) );
  XOR3X2_RVT S2_10_21 ( .A1(ab_10__21_), .A2(CARRYB_9__21_), .A3(SUMB_9__22_), 
        .Y(SUMB_10__21_) );
  XOR3X1_RVT S2_19_12 ( .A1(ab_19__12_), .A2(CARRYB_18__12_), .A3(SUMB_18__13_), .Y(SUMB_19__12_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  AND2X1_RVT U2 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(CARRYB_1__22_) );
  AND2X2_RVT U3 ( .A1(n496), .A2(B[19]), .Y(ab_0__19_) );
  XOR2X1_RVT U4 ( .A1(n348), .A2(n284), .Y(SUMB_1__25_) );
  XOR3X2_RVT U5 ( .A1(ab_2__21_), .A2(CARRYB_1__21_), .A3(SUMB_1__22_), .Y(n3)
         );
  XOR2X2_RVT U6 ( .A1(n236), .A2(n28), .Y(SUMB_1__21_) );
  IBUFFX2_RVT U7 ( .A(n459), .Y(n4) );
  INVX1_RVT U8 ( .A(n4), .Y(n5) );
  AND2X1_RVT U9 ( .A1(n53), .A2(B[23]), .Y(ab_1__23_) );
  NBUFFX2_RVT U10 ( .A(n339), .Y(n6) );
  AND2X4_RVT U11 ( .A1(A[1]), .A2(B[22]), .Y(ab_1__22_) );
  AND2X4_RVT U12 ( .A1(n497), .A2(B[24]), .Y(n250) );
  AND2X4_RVT U13 ( .A1(n53), .A2(B[10]), .Y(ab_1__10_) );
  AND2X1_RVT U14 ( .A1(ab_1__20_), .A2(n138), .Y(n7) );
  NBUFFX2_RVT U15 ( .A(SUMB_25__4_), .Y(n8) );
  NBUFFX2_RVT U16 ( .A(CARRYB_9__18_), .Y(n9) );
  NAND3X0_RVT U17 ( .A1(n323), .A2(n324), .A3(n322), .Y(n10) );
  XOR3X2_RVT U18 ( .A1(SUMB_10__7_), .A2(ab_11__6_), .A3(CARRYB_10__6_), .Y(
        SUMB_11__6_) );
  NAND2X0_RVT U19 ( .A1(SUMB_10__7_), .A2(CARRYB_10__6_), .Y(n11) );
  NAND2X0_RVT U20 ( .A1(ab_11__6_), .A2(CARRYB_10__6_), .Y(n12) );
  NAND2X0_RVT U21 ( .A1(ab_11__6_), .A2(SUMB_10__7_), .Y(n13) );
  NAND3X0_RVT U22 ( .A1(n13), .A2(n12), .A3(n11), .Y(CARRYB_11__6_) );
  AND2X1_RVT U23 ( .A1(n463), .A2(A[1]), .Y(ab_1__20_) );
  AND2X1_RVT U24 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(n14) );
  AND2X4_RVT U25 ( .A1(n53), .A2(B[16]), .Y(ab_1__16_) );
  AND2X4_RVT U26 ( .A1(n250), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X4_RVT U27 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X4_RVT U28 ( .A1(n53), .A2(B[16]), .Y(n327) );
  AND2X4_RVT U29 ( .A1(n54), .A2(B[15]), .Y(ab_1__15_) );
  AND2X4_RVT U30 ( .A1(n53), .A2(B[0]), .Y(ab_1__0_) );
  AND2X4_RVT U31 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  XOR2X1_RVT U32 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(SUMB_1__13_) );
  AND2X4_RVT U33 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  NBUFFX2_RVT U34 ( .A(n340), .Y(n15) );
  XOR2X2_RVT U35 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  NOR2X4_RVT U36 ( .A1(n28), .A2(n236), .Y(CARRYB_1__21_) );
  XOR3X1_RVT U37 ( .A1(CARRYB_14__1_), .A2(ab_15__1_), .A3(SUMB_14__2_), .Y(
        SUMB_15__1_) );
  NAND2X0_RVT U38 ( .A1(SUMB_14__2_), .A2(CARRYB_14__1_), .Y(n16) );
  NAND2X0_RVT U39 ( .A1(ab_15__1_), .A2(CARRYB_14__1_), .Y(n17) );
  NAND2X0_RVT U40 ( .A1(ab_15__1_), .A2(SUMB_14__2_), .Y(n18) );
  NAND3X0_RVT U41 ( .A1(n18), .A2(n17), .A3(n16), .Y(CARRYB_15__1_) );
  XOR3X2_RVT U42 ( .A1(SUMB_15__2_), .A2(ab_16__1_), .A3(CARRYB_15__1_), .Y(
        SUMB_16__1_) );
  NAND2X0_RVT U43 ( .A1(CARRYB_15__1_), .A2(SUMB_15__2_), .Y(n19) );
  NAND2X0_RVT U44 ( .A1(ab_16__1_), .A2(SUMB_15__2_), .Y(n20) );
  NAND2X0_RVT U45 ( .A1(ab_16__1_), .A2(CARRYB_15__1_), .Y(n21) );
  NAND3X0_RVT U46 ( .A1(n21), .A2(n20), .A3(n19), .Y(CARRYB_16__1_) );
  XOR2X2_RVT U47 ( .A1(n23), .A2(n22), .Y(SUMB_1__19_) );
  NAND2X0_RVT U48 ( .A1(n463), .A2(n496), .Y(n22) );
  NAND2X0_RVT U49 ( .A1(B[19]), .A2(n497), .Y(n23) );
  NAND3X2_RVT U50 ( .A1(n292), .A2(n294), .A3(n293), .Y(CARRYB_7__13_) );
  DELLN3X2_RVT U51 ( .A(n456), .Y(n24) );
  AND2X4_RVT U52 ( .A1(n53), .A2(B[12]), .Y(ab_1__12_) );
  AND2X4_RVT U53 ( .A1(n54), .A2(B[29]), .Y(ab_1__29_) );
  AND2X4_RVT U54 ( .A1(n54), .A2(n483), .Y(ab_1__1_) );
  AND2X1_RVT U55 ( .A1(n325), .A2(B[11]), .Y(ab_0__11_) );
  NBUFFX2_RVT U56 ( .A(B[21]), .Y(n148) );
  XOR3X2_RVT U57 ( .A1(CARRYB_3__6_), .A2(ab_4__6_), .A3(SUMB_3__7_), .Y(
        SUMB_4__6_) );
  NAND2X0_RVT U58 ( .A1(SUMB_3__7_), .A2(CARRYB_3__6_), .Y(n25) );
  NAND2X0_RVT U59 ( .A1(ab_4__6_), .A2(CARRYB_3__6_), .Y(n26) );
  NAND2X0_RVT U60 ( .A1(ab_4__6_), .A2(SUMB_3__7_), .Y(n27) );
  NAND3X0_RVT U61 ( .A1(n27), .A2(n26), .A3(n25), .Y(CARRYB_4__6_) );
  AND2X4_RVT U62 ( .A1(n503), .A2(n493), .Y(ab_4__6_) );
  NBUFFX2_RVT U63 ( .A(B[19]), .Y(n462) );
  AND2X1_RVT U64 ( .A1(n508), .A2(n462), .Y(ab_7__19_) );
  OR3X1_RVT U65 ( .A1(n91), .A2(n92), .A3(n93), .Y(CARRYB_5__15_) );
  NAND3X1_RVT U66 ( .A1(n287), .A2(n286), .A3(n285), .Y(CARRYB_8__11_) );
  NAND3X2_RVT U67 ( .A1(n341), .A2(n15), .A3(n6), .Y(n219) );
  NAND3X2_RVT U68 ( .A1(n15), .A2(n341), .A3(n6), .Y(n29) );
  NAND3X2_RVT U69 ( .A1(n345), .A2(n347), .A3(n346), .Y(n189) );
  AND2X4_RVT U70 ( .A1(n148), .A2(n513), .Y(ab_9__21_) );
  NAND2X0_RVT U71 ( .A1(B[21]), .A2(A[1]), .Y(n28) );
  XOR2X1_RVT U72 ( .A1(CARRYB_17__12_), .A2(ab_18__12_), .Y(n30) );
  XOR2X1_RVT U73 ( .A1(SUMB_17__13_), .A2(n30), .Y(SUMB_18__12_) );
  NAND2X0_RVT U74 ( .A1(CARRYB_17__12_), .A2(SUMB_17__13_), .Y(n31) );
  NAND2X0_RVT U75 ( .A1(ab_18__12_), .A2(SUMB_17__13_), .Y(n32) );
  NAND2X0_RVT U76 ( .A1(ab_18__12_), .A2(CARRYB_17__12_), .Y(n33) );
  NAND3X0_RVT U77 ( .A1(n33), .A2(n32), .A3(n31), .Y(CARRYB_18__12_) );
  NBUFFX2_RVT U78 ( .A(SUMB_4__23_), .Y(n34) );
  XOR3X2_RVT U79 ( .A1(SUMB_2__17_), .A2(ab_3__16_), .A3(CARRYB_2__16_), .Y(
        SUMB_3__16_) );
  NAND2X0_RVT U80 ( .A1(CARRYB_2__16_), .A2(SUMB_2__17_), .Y(n35) );
  NAND2X0_RVT U81 ( .A1(ab_3__16_), .A2(SUMB_2__17_), .Y(n36) );
  NAND2X0_RVT U82 ( .A1(ab_3__16_), .A2(CARRYB_2__16_), .Y(n37) );
  NAND3X0_RVT U83 ( .A1(n37), .A2(n36), .A3(n35), .Y(CARRYB_3__16_) );
  AND2X1_RVT U84 ( .A1(n325), .A2(B[17]), .Y(ab_0__17_) );
  XOR2X2_RVT U85 ( .A1(ab_6__21_), .A2(CARRYB_5__21_), .Y(n194) );
  NAND3X2_RVT U86 ( .A1(n206), .A2(n205), .A3(n204), .Y(CARRYB_5__21_) );
  NAND3X2_RVT U87 ( .A1(n76), .A2(n75), .A3(n74), .Y(CARRYB_8__2_) );
  XOR3X2_RVT U88 ( .A1(CARRYB_2__21_), .A2(ab_3__21_), .A3(n131), .Y(n38) );
  DELLN2X2_RVT U89 ( .A(n494), .Y(n39) );
  XOR3X2_RVT U90 ( .A1(SUMB_7__5_), .A2(ab_8__4_), .A3(CARRYB_7__4_), .Y(
        SUMB_8__4_) );
  NAND2X0_RVT U91 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Y(n40) );
  NAND2X0_RVT U92 ( .A1(ab_8__4_), .A2(CARRYB_7__4_), .Y(n41) );
  NAND2X0_RVT U93 ( .A1(ab_8__4_), .A2(SUMB_7__5_), .Y(n42) );
  NAND3X0_RVT U94 ( .A1(n42), .A2(n41), .A3(n40), .Y(CARRYB_8__4_) );
  XOR3X2_RVT U95 ( .A1(SUMB_12__4_), .A2(ab_13__3_), .A3(CARRYB_12__3_), .Y(
        SUMB_13__3_) );
  NAND2X0_RVT U96 ( .A1(CARRYB_12__3_), .A2(SUMB_12__4_), .Y(n43) );
  NAND2X0_RVT U97 ( .A1(ab_13__3_), .A2(SUMB_12__4_), .Y(n44) );
  NAND2X0_RVT U98 ( .A1(ab_13__3_), .A2(CARRYB_12__3_), .Y(n45) );
  NAND3X0_RVT U99 ( .A1(n45), .A2(n44), .A3(n43), .Y(CARRYB_13__3_) );
  NAND3X1_RVT U100 ( .A1(n52), .A2(n51), .A3(n50), .Y(CARRYB_7__4_) );
  AND2X4_RVT U101 ( .A1(A[5]), .A2(n148), .Y(ab_5__21_) );
  XOR2X2_RVT U102 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  NBUFFX2_RVT U103 ( .A(SUMB_7__18_), .Y(n46) );
  XOR3X2_RVT U104 ( .A1(CARRYB_11__4_), .A2(ab_12__4_), .A3(SUMB_11__5_), .Y(
        SUMB_12__4_) );
  NAND2X0_RVT U105 ( .A1(SUMB_11__5_), .A2(CARRYB_11__4_), .Y(n47) );
  NAND2X0_RVT U106 ( .A1(ab_12__4_), .A2(CARRYB_11__4_), .Y(n48) );
  NAND2X0_RVT U107 ( .A1(ab_12__4_), .A2(SUMB_11__5_), .Y(n49) );
  NAND3X0_RVT U108 ( .A1(n49), .A2(n48), .A3(n47), .Y(CARRYB_12__4_) );
  XOR3X2_RVT U109 ( .A1(CARRYB_6__4_), .A2(ab_7__4_), .A3(SUMB_6__5_), .Y(
        SUMB_7__4_) );
  NAND2X0_RVT U110 ( .A1(SUMB_6__5_), .A2(CARRYB_6__4_), .Y(n50) );
  NAND2X0_RVT U111 ( .A1(ab_7__4_), .A2(CARRYB_6__4_), .Y(n51) );
  NAND2X0_RVT U112 ( .A1(ab_7__4_), .A2(SUMB_6__5_), .Y(n52) );
  NBUFFX2_RVT U113 ( .A(B[22]), .Y(n464) );
  NBUFFX2_RVT U114 ( .A(A[1]), .Y(n53) );
  NBUFFX2_RVT U115 ( .A(A[1]), .Y(n54) );
  INVX0_RVT U116 ( .A(n493), .Y(n55) );
  IBUFFX8_RVT U117 ( .A(n55), .Y(n56) );
  AND2X4_RVT U118 ( .A1(n56), .A2(n513), .Y(ab_9__6_) );
  NBUFFX2_RVT U119 ( .A(A[0]), .Y(n57) );
  NAND3X0_RVT U120 ( .A1(n106), .A2(n105), .A3(n104), .Y(n58) );
  NAND3X0_RVT U121 ( .A1(n106), .A2(n105), .A3(n104), .Y(n59) );
  XOR3X2_RVT U122 ( .A1(CARRYB_10__2_), .A2(ab_11__2_), .A3(SUMB_10__3_), .Y(
        SUMB_11__2_) );
  NAND2X0_RVT U123 ( .A1(SUMB_10__3_), .A2(CARRYB_10__2_), .Y(n60) );
  NAND2X0_RVT U124 ( .A1(ab_11__2_), .A2(CARRYB_10__2_), .Y(n61) );
  NAND2X0_RVT U125 ( .A1(ab_11__2_), .A2(SUMB_10__3_), .Y(n62) );
  NAND3X0_RVT U126 ( .A1(n62), .A2(n61), .A3(n60), .Y(CARRYB_11__2_) );
  NAND3X0_RVT U127 ( .A1(n385), .A2(n386), .A3(n384), .Y(CARRYB_3__20_) );
  AND2X1_RVT U128 ( .A1(n508), .A2(n220), .Y(ab_7__18_) );
  NAND3X0_RVT U129 ( .A1(n365), .A2(n364), .A3(n363), .Y(CARRYB_6__18_) );
  XOR2X1_RVT U130 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(SUMB_1__12_) );
  NAND3X0_RVT U131 ( .A1(n126), .A2(n127), .A3(n125), .Y(CARRYB_6__3_) );
  AND2X1_RVT U132 ( .A1(n167), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U133 ( .A1(ab_1__28_), .A2(n406), .Y(CARRYB_1__28_) );
  NAND2X0_RVT U134 ( .A1(ab_3__14_), .A2(CARRYB_2__14_), .Y(n103) );
  AND2X1_RVT U135 ( .A1(n501), .A2(B[24]), .Y(ab_3__24_) );
  NAND3X0_RVT U136 ( .A1(n121), .A2(n120), .A3(n119), .Y(CARRYB_4__20_) );
  NAND3X0_RVT U137 ( .A1(n109), .A2(n108), .A3(n107), .Y(CARRYB_7__18_) );
  NAND2X0_RVT U138 ( .A1(ab_7__18_), .A2(CARRYB_6__18_), .Y(n109) );
  NAND3X1_RVT U139 ( .A1(n359), .A2(n358), .A3(n357), .Y(CARRYB_10__18_) );
  AND2X1_RVT U140 ( .A1(n143), .A2(n512), .Y(ab_9__16_) );
  NAND3X0_RVT U141 ( .A1(n100), .A2(n99), .A3(n98), .Y(CARRYB_9__17_) );
  NAND2X0_RVT U142 ( .A1(ab_3__10_), .A2(CARRYB_2__10_), .Y(n70) );
  AND2X1_RVT U143 ( .A1(n501), .A2(n495), .Y(ab_3__9_) );
  XOR2X1_RVT U144 ( .A1(n162), .A2(SUMB_12__16_), .Y(SUMB_13__15_) );
  NAND3X0_RVT U145 ( .A1(n223), .A2(n222), .A3(n221), .Y(CARRYB_26__3_) );
  NAND2X0_RVT U146 ( .A1(ab_8__2_), .A2(CARRYB_7__2_), .Y(n76) );
  AND2X1_RVT U147 ( .A1(n484), .A2(n512), .Y(ab_9__1_) );
  NAND3X0_RVT U148 ( .A1(n83), .A2(n82), .A3(n81), .Y(CARRYB_12__1_) );
  NAND2X0_RVT U149 ( .A1(ab_27__0_), .A2(CARRYB_26__0_), .Y(n124) );
  XOR3X2_RVT U150 ( .A1(SUMB_6__4_), .A2(ab_7__3_), .A3(CARRYB_6__3_), .Y(
        SUMB_7__3_) );
  NAND2X0_RVT U151 ( .A1(CARRYB_6__3_), .A2(SUMB_6__4_), .Y(n63) );
  NAND2X0_RVT U152 ( .A1(ab_7__3_), .A2(SUMB_6__4_), .Y(n64) );
  NAND2X0_RVT U153 ( .A1(ab_7__3_), .A2(CARRYB_6__3_), .Y(n65) );
  NAND3X0_RVT U154 ( .A1(n65), .A2(n64), .A3(n63), .Y(CARRYB_7__3_) );
  XOR2X2_RVT U155 ( .A1(CARRYB_1__28_), .A2(ab_2__28_), .Y(n66) );
  XOR2X2_RVT U156 ( .A1(SUMB_1__29_), .A2(n66), .Y(SUMB_2__28_) );
  XOR2X1_RVT U157 ( .A1(CARRYB_9__20_), .A2(ab_10__20_), .Y(n67) );
  XOR2X2_RVT U158 ( .A1(SUMB_9__21_), .A2(n67), .Y(SUMB_10__20_) );
  XOR2X2_RVT U159 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(SUMB_1__17_) );
  XOR3X2_RVT U160 ( .A1(SUMB_2__11_), .A2(ab_3__10_), .A3(CARRYB_2__10_), .Y(
        SUMB_3__10_) );
  NAND2X0_RVT U161 ( .A1(CARRYB_2__10_), .A2(SUMB_2__11_), .Y(n68) );
  NAND2X0_RVT U162 ( .A1(ab_3__10_), .A2(SUMB_2__11_), .Y(n69) );
  NAND3X0_RVT U163 ( .A1(n70), .A2(n69), .A3(n68), .Y(CARRYB_3__10_) );
  XOR3X2_RVT U164 ( .A1(CARRYB_8__8_), .A2(ab_9__8_), .A3(SUMB_8__9_), .Y(
        SUMB_9__8_) );
  NAND2X0_RVT U165 ( .A1(SUMB_8__9_), .A2(CARRYB_8__8_), .Y(n71) );
  NAND2X0_RVT U166 ( .A1(ab_9__8_), .A2(CARRYB_8__8_), .Y(n72) );
  NAND2X0_RVT U167 ( .A1(ab_9__8_), .A2(SUMB_8__9_), .Y(n73) );
  NAND3X0_RVT U168 ( .A1(n73), .A2(n72), .A3(n71), .Y(CARRYB_9__8_) );
  NAND2X0_RVT U169 ( .A1(ab_5__9_), .A2(CARRYB_4__9_), .Y(n137) );
  XOR3X2_RVT U170 ( .A1(SUMB_7__3_), .A2(ab_8__2_), .A3(CARRYB_7__2_), .Y(
        SUMB_8__2_) );
  NAND2X0_RVT U171 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Y(n74) );
  NAND2X0_RVT U172 ( .A1(ab_8__2_), .A2(SUMB_7__3_), .Y(n75) );
  XOR3X2_RVT U173 ( .A1(SUMB_8__3_), .A2(ab_9__2_), .A3(CARRYB_8__2_), .Y(
        SUMB_9__2_) );
  NAND2X0_RVT U174 ( .A1(CARRYB_8__2_), .A2(SUMB_8__3_), .Y(n77) );
  NAND2X0_RVT U175 ( .A1(ab_9__2_), .A2(SUMB_8__3_), .Y(n78) );
  NAND2X0_RVT U176 ( .A1(ab_9__2_), .A2(CARRYB_8__2_), .Y(n79) );
  NAND3X0_RVT U177 ( .A1(n79), .A2(n78), .A3(n77), .Y(CARRYB_9__2_) );
  AND2X4_RVT U178 ( .A1(n485), .A2(n513), .Y(ab_9__2_) );
  NAND3X0_RVT U179 ( .A1(n329), .A2(n330), .A3(n328), .Y(n80) );
  AND2X4_RVT U180 ( .A1(n381), .A2(n482), .Y(PRODUCT_0_) );
  XOR2X1_RVT U181 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U182 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR3X2_RVT U183 ( .A1(CARRYB_11__1_), .A2(ab_12__1_), .A3(SUMB_11__2_), .Y(
        SUMB_12__1_) );
  NAND2X0_RVT U184 ( .A1(SUMB_11__2_), .A2(CARRYB_11__1_), .Y(n81) );
  NAND2X0_RVT U185 ( .A1(ab_12__1_), .A2(CARRYB_11__1_), .Y(n82) );
  NAND2X0_RVT U186 ( .A1(ab_12__1_), .A2(SUMB_11__2_), .Y(n83) );
  XOR3X2_RVT U187 ( .A1(SUMB_12__2_), .A2(ab_13__1_), .A3(CARRYB_12__1_), .Y(
        SUMB_13__1_) );
  NAND2X0_RVT U188 ( .A1(CARRYB_12__1_), .A2(SUMB_12__2_), .Y(n84) );
  NAND2X0_RVT U189 ( .A1(ab_13__1_), .A2(SUMB_12__2_), .Y(n85) );
  NAND2X0_RVT U190 ( .A1(ab_13__1_), .A2(CARRYB_12__1_), .Y(n86) );
  NAND3X0_RVT U191 ( .A1(n86), .A2(n85), .A3(n84), .Y(CARRYB_13__1_) );
  XOR3X2_RVT U192 ( .A1(CARRYB_8__1_), .A2(ab_9__1_), .A3(SUMB_8__2_), .Y(
        SUMB_9__1_) );
  NAND2X0_RVT U193 ( .A1(SUMB_8__2_), .A2(CARRYB_8__1_), .Y(n87) );
  NAND2X0_RVT U194 ( .A1(ab_9__1_), .A2(CARRYB_8__1_), .Y(n88) );
  NAND2X0_RVT U195 ( .A1(ab_9__1_), .A2(SUMB_8__2_), .Y(n89) );
  NAND3X0_RVT U196 ( .A1(n89), .A2(n88), .A3(n87), .Y(CARRYB_9__1_) );
  NBUFFX2_RVT U197 ( .A(SUMB_4__21_), .Y(n90) );
  AND2X1_RVT U198 ( .A1(ab_5__15_), .A2(CARRYB_4__15_), .Y(n91) );
  AND2X1_RVT U199 ( .A1(ab_5__15_), .A2(SUMB_4__16_), .Y(n92) );
  AND2X1_RVT U200 ( .A1(SUMB_4__16_), .A2(CARRYB_4__15_), .Y(n93) );
  IBUFFX2_RVT U201 ( .A(n463), .Y(n276) );
  XOR3X2_RVT U202 ( .A1(n94), .A2(n95), .A3(n96), .Y(n114) );
  NAND2X0_RVT U203 ( .A1(A[28]), .A2(n487), .Y(n94) );
  AND3X1_RVT U204 ( .A1(n428), .A2(n427), .A3(n426), .Y(n95) );
  XNOR3X2_RVT U205 ( .A1(ab_27__4_), .A2(CARRYB_26__4_), .A3(SUMB_26__5_), .Y(
        n96) );
  NAND3X0_RVT U206 ( .A1(n154), .A2(n153), .A3(n152), .Y(n97) );
  XOR3X2_RVT U207 ( .A1(CARRYB_8__17_), .A2(ab_9__17_), .A3(SUMB_8__18_), .Y(
        SUMB_9__17_) );
  NAND2X0_RVT U208 ( .A1(SUMB_8__18_), .A2(n59), .Y(n98) );
  NAND2X0_RVT U209 ( .A1(ab_9__17_), .A2(n58), .Y(n99) );
  NAND2X0_RVT U210 ( .A1(ab_9__17_), .A2(SUMB_8__18_), .Y(n100) );
  XOR3X2_RVT U211 ( .A1(CARRYB_2__14_), .A2(ab_3__14_), .A3(SUMB_2__15_), .Y(
        SUMB_3__14_) );
  NAND2X0_RVT U212 ( .A1(CARRYB_2__14_), .A2(SUMB_2__15_), .Y(n101) );
  NAND2X0_RVT U213 ( .A1(ab_3__14_), .A2(SUMB_2__15_), .Y(n102) );
  NAND3X0_RVT U214 ( .A1(n102), .A2(n103), .A3(n101), .Y(CARRYB_3__14_) );
  XOR3X2_RVT U215 ( .A1(CARRYB_7__17_), .A2(ab_8__17_), .A3(n46), .Y(
        SUMB_8__17_) );
  NAND2X0_RVT U216 ( .A1(CARRYB_7__17_), .A2(SUMB_7__18_), .Y(n104) );
  NAND2X0_RVT U217 ( .A1(ab_8__17_), .A2(SUMB_7__18_), .Y(n105) );
  NAND2X0_RVT U218 ( .A1(ab_8__17_), .A2(CARRYB_7__17_), .Y(n106) );
  NAND3X0_RVT U219 ( .A1(n105), .A2(n106), .A3(n104), .Y(CARRYB_8__17_) );
  XOR3X2_RVT U220 ( .A1(CARRYB_6__18_), .A2(ab_7__18_), .A3(SUMB_6__19_), .Y(
        SUMB_7__18_) );
  NAND2X0_RVT U221 ( .A1(CARRYB_6__18_), .A2(SUMB_6__19_), .Y(n107) );
  NAND2X0_RVT U222 ( .A1(ab_7__18_), .A2(SUMB_6__19_), .Y(n108) );
  NAND2X0_RVT U223 ( .A1(ab_8__18_), .A2(CARRYB_7__18_), .Y(n134) );
  XOR2X2_RVT U224 ( .A1(n198), .A2(n178), .Y(SUMB_1__20_) );
  NBUFFX2_RVT U225 ( .A(CARRYB_28__1_), .Y(n110) );
  NAND3X0_RVT U226 ( .A1(n434), .A2(n433), .A3(n432), .Y(n111) );
  NAND3X0_RVT U227 ( .A1(n434), .A2(n433), .A3(n432), .Y(CARRYB_27__2_) );
  XOR3X2_RVT U228 ( .A1(n112), .A2(n113), .A3(n114), .Y(n139) );
  NAND2X0_RVT U229 ( .A1(A[29]), .A2(n485), .Y(n112) );
  AND3X1_RVT U230 ( .A1(n440), .A2(n439), .A3(n438), .Y(n113) );
  AND2X1_RVT U231 ( .A1(n498), .A2(n161), .Y(n115) );
  XOR3X2_RVT U232 ( .A1(CARRYB_6__19_), .A2(ab_7__19_), .A3(SUMB_6__20_), .Y(
        SUMB_7__19_) );
  NAND2X0_RVT U233 ( .A1(SUMB_6__20_), .A2(CARRYB_6__19_), .Y(n116) );
  NAND2X0_RVT U234 ( .A1(ab_7__19_), .A2(CARRYB_6__19_), .Y(n117) );
  NAND2X0_RVT U235 ( .A1(ab_7__19_), .A2(SUMB_6__20_), .Y(n118) );
  NAND3X0_RVT U236 ( .A1(n118), .A2(n117), .A3(n116), .Y(CARRYB_7__19_) );
  XOR3X2_RVT U237 ( .A1(SUMB_3__21_), .A2(ab_4__20_), .A3(CARRYB_3__20_), .Y(
        SUMB_4__20_) );
  NAND2X0_RVT U238 ( .A1(CARRYB_3__20_), .A2(n38), .Y(n119) );
  NAND2X0_RVT U239 ( .A1(ab_4__20_), .A2(n38), .Y(n120) );
  NAND2X0_RVT U240 ( .A1(ab_4__20_), .A2(CARRYB_3__20_), .Y(n121) );
  XOR3X2_RVT U241 ( .A1(SUMB_26__1_), .A2(ab_27__0_), .A3(CARRYB_26__0_), .Y(
        PRODUCT_27_) );
  NAND2X0_RVT U242 ( .A1(CARRYB_26__0_), .A2(SUMB_26__1_), .Y(n122) );
  NAND2X0_RVT U243 ( .A1(ab_27__0_), .A2(SUMB_26__1_), .Y(n123) );
  NAND3X0_RVT U244 ( .A1(n124), .A2(n123), .A3(n122), .Y(CARRYB_27__0_) );
  XOR3X2_RVT U245 ( .A1(n97), .A2(ab_6__3_), .A3(SUMB_5__4_), .Y(SUMB_6__3_)
         );
  NAND2X0_RVT U246 ( .A1(SUMB_5__4_), .A2(CARRYB_5__3_), .Y(n125) );
  NAND2X0_RVT U247 ( .A1(ab_6__3_), .A2(CARRYB_5__3_), .Y(n126) );
  NAND2X0_RVT U248 ( .A1(ab_6__3_), .A2(SUMB_5__4_), .Y(n127) );
  XOR3X1_RVT U249 ( .A1(SUMB_20__1_), .A2(ab_21__0_), .A3(CARRYB_20__0_), .Y(
        PRODUCT_21_) );
  NAND2X0_RVT U250 ( .A1(CARRYB_20__0_), .A2(SUMB_20__1_), .Y(n128) );
  NAND2X0_RVT U251 ( .A1(ab_21__0_), .A2(SUMB_20__1_), .Y(n129) );
  NAND2X0_RVT U252 ( .A1(ab_21__0_), .A2(CARRYB_20__0_), .Y(n130) );
  NAND3X0_RVT U253 ( .A1(n130), .A2(n129), .A3(n128), .Y(CARRYB_21__0_) );
  XOR3X2_RVT U254 ( .A1(ab_2__22_), .A2(CARRYB_1__22_), .A3(SUMB_1__23_), .Y(
        n131) );
  AND2X1_RVT U255 ( .A1(n510), .A2(n220), .Y(ab_8__18_) );
  XOR3X2_RVT U256 ( .A1(SUMB_7__19_), .A2(ab_8__18_), .A3(CARRYB_7__18_), .Y(
        SUMB_8__18_) );
  NAND2X0_RVT U257 ( .A1(CARRYB_7__18_), .A2(SUMB_7__19_), .Y(n132) );
  NAND2X0_RVT U258 ( .A1(ab_8__18_), .A2(SUMB_7__19_), .Y(n133) );
  NAND3X0_RVT U259 ( .A1(n134), .A2(n133), .A3(n132), .Y(CARRYB_8__18_) );
  XOR2X2_RVT U260 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR3X2_RVT U261 ( .A1(CARRYB_4__9_), .A2(ab_5__9_), .A3(SUMB_4__10_), .Y(
        SUMB_5__9_) );
  NAND2X0_RVT U262 ( .A1(CARRYB_4__9_), .A2(SUMB_4__10_), .Y(n135) );
  NAND2X0_RVT U263 ( .A1(ab_5__9_), .A2(SUMB_4__10_), .Y(n136) );
  NAND3X0_RVT U264 ( .A1(n137), .A2(n136), .A3(n135), .Y(CARRYB_5__9_) );
  AND2X4_RVT U265 ( .A1(n505), .A2(n238), .Y(ab_5__9_) );
  AND2X1_RVT U266 ( .A1(n496), .A2(n463), .Y(ab_0__20_) );
  INVX0_RVT U267 ( .A(n178), .Y(n138) );
  XOR3X2_RVT U268 ( .A1(n350), .A2(n349), .A3(n139), .Y(n343) );
  XOR3X2_RVT U269 ( .A1(SUMB_4__21_), .A2(ab_5__20_), .A3(CARRYB_4__20_), .Y(
        SUMB_5__20_) );
  NAND2X0_RVT U270 ( .A1(CARRYB_4__20_), .A2(n90), .Y(n140) );
  NAND2X0_RVT U271 ( .A1(ab_5__20_), .A2(n90), .Y(n141) );
  NAND2X0_RVT U272 ( .A1(ab_5__20_), .A2(CARRYB_4__20_), .Y(n142) );
  NAND3X0_RVT U273 ( .A1(n142), .A2(n141), .A3(n140), .Y(CARRYB_5__20_) );
  NBUFFX2_RVT U274 ( .A(B[16]), .Y(n143) );
  NAND3X0_RVT U275 ( .A1(n313), .A2(n314), .A3(n312), .Y(n144) );
  XOR3X2_RVT U276 ( .A1(SUMB_5__21_), .A2(ab_6__20_), .A3(CARRYB_5__20_), .Y(
        SUMB_6__20_) );
  NAND2X0_RVT U277 ( .A1(CARRYB_5__20_), .A2(SUMB_5__21_), .Y(n145) );
  NAND2X0_RVT U278 ( .A1(ab_6__20_), .A2(SUMB_5__21_), .Y(n146) );
  NAND2X0_RVT U279 ( .A1(ab_6__20_), .A2(CARRYB_5__20_), .Y(n147) );
  NAND3X0_RVT U280 ( .A1(n147), .A2(n146), .A3(n145), .Y(CARRYB_6__20_) );
  AND2X1_RVT U281 ( .A1(n507), .A2(n148), .Y(ab_6__21_) );
  XOR3X2_RVT U282 ( .A1(CARRYB_3__5_), .A2(ab_4__5_), .A3(SUMB_3__6_), .Y(
        SUMB_4__5_) );
  NAND2X0_RVT U283 ( .A1(CARRYB_3__5_), .A2(SUMB_3__6_), .Y(n149) );
  NAND2X0_RVT U284 ( .A1(ab_4__5_), .A2(CARRYB_3__5_), .Y(n150) );
  NAND2X0_RVT U285 ( .A1(ab_4__5_), .A2(SUMB_3__6_), .Y(n151) );
  NAND3X0_RVT U286 ( .A1(n151), .A2(n150), .A3(n149), .Y(CARRYB_4__5_) );
  XOR3X2_RVT U287 ( .A1(SUMB_4__4_), .A2(ab_5__3_), .A3(CARRYB_4__3_), .Y(
        SUMB_5__3_) );
  NAND2X0_RVT U288 ( .A1(CARRYB_4__3_), .A2(SUMB_4__4_), .Y(n152) );
  NAND2X0_RVT U289 ( .A1(ab_5__3_), .A2(SUMB_4__4_), .Y(n153) );
  NAND2X0_RVT U290 ( .A1(ab_5__3_), .A2(CARRYB_4__3_), .Y(n154) );
  NAND3X0_RVT U291 ( .A1(n154), .A2(n153), .A3(n152), .Y(CARRYB_5__3_) );
  NBUFFX2_RVT U292 ( .A(CARRYB_29__0_), .Y(n155) );
  XOR3X2_RVT U293 ( .A1(CARRYB_2__22_), .A2(ab_3__22_), .A3(SUMB_2__23_), .Y(
        SUMB_3__22_) );
  NAND2X0_RVT U294 ( .A1(SUMB_2__23_), .A2(CARRYB_2__22_), .Y(n156) );
  NAND2X0_RVT U295 ( .A1(ab_3__22_), .A2(CARRYB_2__22_), .Y(n157) );
  NAND2X0_RVT U296 ( .A1(ab_3__22_), .A2(SUMB_2__23_), .Y(n158) );
  NAND3X0_RVT U297 ( .A1(n158), .A2(n157), .A3(n156), .Y(CARRYB_3__22_) );
  NAND3X0_RVT U298 ( .A1(n308), .A2(n307), .A3(n306), .Y(n159) );
  NAND3X0_RVT U299 ( .A1(n308), .A2(n307), .A3(n306), .Y(n160) );
  NAND2X0_RVT U300 ( .A1(ab_2__27_), .A2(CARRYB_1__27_), .Y(n275) );
  AND2X1_RVT U301 ( .A1(n381), .A2(B[27]), .Y(ab_0__27_) );
  NAND3X0_RVT U302 ( .A1(n399), .A2(n398), .A3(n397), .Y(CARRYB_2__26_) );
  NAND3X0_RVT U303 ( .A1(n321), .A2(n320), .A3(n319), .Y(CARRYB_7__11_) );
  NAND3X0_RVT U304 ( .A1(n437), .A2(n436), .A3(n435), .Y(CARRYB_7__22_) );
  NAND3X0_RVT U305 ( .A1(n418), .A2(n417), .A3(n416), .Y(CARRYB_12__17_) );
  AND2X1_RVT U306 ( .A1(n248), .A2(n490), .Y(ab_2__4_) );
  AND2X1_RVT U307 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U308 ( .A1(n248), .A2(n485), .Y(ab_2__2_) );
  AND2X1_RVT U309 ( .A1(n248), .A2(n488), .Y(ab_2__3_) );
  AND2X1_RVT U310 ( .A1(n501), .A2(n299), .Y(ab_3__23_) );
  INVX1_RVT U311 ( .A(n331), .Y(n332) );
  NAND3X0_RVT U312 ( .A1(n393), .A2(n392), .A3(n391), .Y(CARRYB_4__24_) );
  AND2X1_RVT U313 ( .A1(n325), .A2(B[13]), .Y(ab_0__13_) );
  AND2X1_RVT U314 ( .A1(n507), .A2(n457), .Y(ab_6__12_) );
  NAND3X0_RVT U315 ( .A1(n380), .A2(n379), .A3(n378), .Y(CARRYB_6__22_) );
  NAND3X0_RVT U316 ( .A1(n259), .A2(n258), .A3(n257), .Y(CARRYB_8__20_) );
  AND2X1_RVT U317 ( .A1(n220), .A2(n512), .Y(ab_9__18_) );
  AND2X1_RVT U318 ( .A1(n224), .A2(n512), .Y(ab_9__17_) );
  XOR2X1_RVT U319 ( .A1(CARRYB_12__15_), .A2(ab_13__15_), .Y(n162) );
  NAND3X0_RVT U320 ( .A1(n421), .A2(n420), .A3(n419), .Y(CARRYB_15__14_) );
  NAND3X0_RVT U321 ( .A1(n405), .A2(n404), .A3(n403), .Y(CARRYB_25__4_) );
  AND2X1_RVT U322 ( .A1(n501), .A2(n488), .Y(ab_3__3_) );
  NAND3X0_RVT U323 ( .A1(n402), .A2(n401), .A3(n400), .Y(CARRYB_26__2_) );
  NAND3X0_RVT U324 ( .A1(n184), .A2(n183), .A3(n182), .Y(CARRYB_4__1_) );
  AND2X1_RVT U325 ( .A1(n167), .A2(n484), .Y(ab_0__1_) );
  AND2X1_RVT U326 ( .A1(n501), .A2(n481), .Y(ab_3__0_) );
  NBUFFX2_RVT U327 ( .A(B[7]), .Y(n161) );
  NAND2X0_RVT U328 ( .A1(CARRYB_12__15_), .A2(SUMB_12__16_), .Y(n163) );
  NAND2X0_RVT U329 ( .A1(ab_13__15_), .A2(SUMB_12__16_), .Y(n164) );
  NAND2X0_RVT U330 ( .A1(ab_13__15_), .A2(CARRYB_12__15_), .Y(n165) );
  NAND3X0_RVT U331 ( .A1(n165), .A2(n164), .A3(n163), .Y(CARRYB_13__15_) );
  XOR3X2_RVT U332 ( .A1(ab_5__22_), .A2(CARRYB_4__22_), .A3(n34), .Y(n166) );
  DELLN3X2_RVT U333 ( .A(n381), .Y(n167) );
  AND2X1_RVT U334 ( .A1(B[25]), .A2(n57), .Y(ab_0__25_) );
  XOR2X2_RVT U335 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  AND2X1_RVT U336 ( .A1(n57), .A2(n492), .Y(ab_0__5_) );
  AND2X1_RVT U337 ( .A1(n498), .A2(n492), .Y(ab_1__5_) );
  AND2X1_RVT U338 ( .A1(B[24]), .A2(n57), .Y(n168) );
  NBUFFX2_RVT U339 ( .A(CARRYB_25__3_), .Y(n169) );
  XOR3X2_RVT U340 ( .A1(CARRYB_26__1_), .A2(ab_27__1_), .A3(SUMB_26__2_), .Y(
        SUMB_27__1_) );
  NAND2X0_RVT U341 ( .A1(SUMB_26__2_), .A2(CARRYB_26__1_), .Y(n170) );
  NAND2X0_RVT U342 ( .A1(ab_27__1_), .A2(CARRYB_26__1_), .Y(n171) );
  NAND2X0_RVT U343 ( .A1(ab_27__1_), .A2(SUMB_26__2_), .Y(n172) );
  NAND3X0_RVT U344 ( .A1(n172), .A2(n171), .A3(n170), .Y(CARRYB_27__1_) );
  NAND3X0_RVT U345 ( .A1(n231), .A2(n232), .A3(n230), .Y(n173) );
  NBUFFX2_RVT U346 ( .A(A[1]), .Y(n497) );
  AND2X1_RVT U347 ( .A1(n503), .A2(n462), .Y(ab_4__19_) );
  AND2X2_RVT U348 ( .A1(n57), .A2(B[29]), .Y(n406) );
  AND2X4_RVT U349 ( .A1(n325), .A2(B[10]), .Y(ab_0__10_) );
  AND2X4_RVT U350 ( .A1(n381), .A2(B[15]), .Y(ab_0__15_) );
  AND2X4_RVT U351 ( .A1(n325), .A2(B[6]), .Y(ab_0__6_) );
  NBUFFX2_RVT U352 ( .A(SUMB_4__8_), .Y(n174) );
  XOR2X1_RVT U353 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  XOR3X2_RVT U354 ( .A1(CARRYB_5__15_), .A2(ab_6__15_), .A3(SUMB_5__16_), .Y(
        SUMB_6__15_) );
  NAND2X0_RVT U355 ( .A1(CARRYB_5__15_), .A2(SUMB_5__16_), .Y(n175) );
  NAND2X0_RVT U356 ( .A1(ab_6__15_), .A2(CARRYB_5__15_), .Y(n176) );
  NAND2X0_RVT U357 ( .A1(ab_6__15_), .A2(SUMB_5__16_), .Y(n177) );
  NAND3X0_RVT U358 ( .A1(n177), .A2(n176), .A3(n175), .Y(CARRYB_6__15_) );
  NAND2X0_RVT U359 ( .A1(B[21]), .A2(A[0]), .Y(n178) );
  XOR3X2_RVT U360 ( .A1(CARRYB_5__1_), .A2(ab_6__1_), .A3(SUMB_5__2_), .Y(
        SUMB_6__1_) );
  NAND2X0_RVT U361 ( .A1(SUMB_5__2_), .A2(CARRYB_5__1_), .Y(n179) );
  NAND2X0_RVT U362 ( .A1(ab_6__1_), .A2(CARRYB_5__1_), .Y(n180) );
  NAND2X0_RVT U363 ( .A1(ab_6__1_), .A2(SUMB_5__2_), .Y(n181) );
  NAND3X0_RVT U364 ( .A1(n181), .A2(n180), .A3(n179), .Y(CARRYB_6__1_) );
  XOR3X2_RVT U365 ( .A1(CARRYB_3__1_), .A2(ab_4__1_), .A3(SUMB_3__2_), .Y(
        SUMB_4__1_) );
  NAND2X0_RVT U366 ( .A1(SUMB_3__2_), .A2(CARRYB_3__1_), .Y(n182) );
  NAND2X0_RVT U367 ( .A1(ab_4__1_), .A2(CARRYB_3__1_), .Y(n183) );
  NAND2X0_RVT U368 ( .A1(ab_4__1_), .A2(SUMB_3__2_), .Y(n184) );
  XOR3X2_RVT U369 ( .A1(CARRYB_4__1_), .A2(ab_5__1_), .A3(SUMB_4__2_), .Y(
        SUMB_5__1_) );
  NAND2X0_RVT U370 ( .A1(SUMB_4__2_), .A2(CARRYB_4__1_), .Y(n185) );
  NAND2X0_RVT U371 ( .A1(ab_5__1_), .A2(CARRYB_4__1_), .Y(n186) );
  NAND2X0_RVT U372 ( .A1(ab_5__1_), .A2(SUMB_4__2_), .Y(n187) );
  NAND3X0_RVT U373 ( .A1(n187), .A2(n186), .A3(n185), .Y(CARRYB_5__1_) );
  NAND3X0_RVT U374 ( .A1(n214), .A2(n215), .A3(n213), .Y(n188) );
  AND2X1_RVT U375 ( .A1(B[23]), .A2(A[0]), .Y(ab_0__23_) );
  NAND3X0_RVT U376 ( .A1(n345), .A2(n346), .A3(n347), .Y(n190) );
  XOR2X2_RVT U377 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR3X2_RVT U378 ( .A1(CARRYB_18__9_), .A2(ab_19__9_), .A3(SUMB_18__10_), .Y(
        SUMB_19__9_) );
  NAND2X0_RVT U379 ( .A1(CARRYB_18__9_), .A2(SUMB_18__10_), .Y(n191) );
  NAND2X0_RVT U380 ( .A1(ab_19__9_), .A2(SUMB_18__10_), .Y(n192) );
  NAND2X0_RVT U381 ( .A1(ab_19__9_), .A2(CARRYB_18__9_), .Y(n193) );
  NAND3X0_RVT U382 ( .A1(n193), .A2(n192), .A3(n191), .Y(CARRYB_19__9_) );
  XOR2X2_RVT U383 ( .A1(n166), .A2(n194), .Y(SUMB_6__21_) );
  NAND2X0_RVT U384 ( .A1(ab_6__21_), .A2(SUMB_5__22_), .Y(n195) );
  NAND2X0_RVT U385 ( .A1(CARRYB_5__21_), .A2(SUMB_5__22_), .Y(n196) );
  NAND2X0_RVT U386 ( .A1(CARRYB_5__21_), .A2(ab_6__21_), .Y(n197) );
  NAND3X2_RVT U387 ( .A1(n197), .A2(n196), .A3(n195), .Y(CARRYB_6__21_) );
  NAND3X0_RVT U388 ( .A1(n362), .A2(n361), .A3(n360), .Y(CARRYB_9__18_) );
  AND2X1_RVT U389 ( .A1(B[24]), .A2(A[0]), .Y(ab_0__24_) );
  NAND2X0_RVT U390 ( .A1(B[20]), .A2(A[1]), .Y(n198) );
  AND2X1_RVT U391 ( .A1(n498), .A2(n487), .Y(ab_1__3_) );
  XOR2X1_RVT U392 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR3X2_RVT U393 ( .A1(ab_8__21_), .A2(CARRYB_7__21_), .A3(SUMB_7__22_), .Y(
        n199) );
  XOR3X2_RVT U394 ( .A1(ab_11__18_), .A2(CARRYB_10__18_), .A3(SUMB_10__19_), 
        .Y(n200) );
  XOR2X1_RVT U395 ( .A1(CARRYB_22__7_), .A2(ab_23__7_), .Y(n201) );
  XOR2X2_RVT U396 ( .A1(SUMB_22__8_), .A2(n201), .Y(SUMB_23__7_) );
  NBUFFX2_RVT U397 ( .A(SUMB_3__22_), .Y(n202) );
  XOR3X2_RVT U398 ( .A1(n169), .A2(ab_26__3_), .A3(n8), .Y(n203) );
  XOR3X2_RVT U399 ( .A1(CARRYB_4__21_), .A2(ab_5__21_), .A3(SUMB_4__22_), .Y(
        SUMB_5__21_) );
  NAND2X0_RVT U400 ( .A1(SUMB_4__22_), .A2(CARRYB_4__21_), .Y(n204) );
  NAND2X0_RVT U401 ( .A1(ab_5__21_), .A2(n188), .Y(n205) );
  NAND2X0_RVT U402 ( .A1(ab_5__21_), .A2(SUMB_4__22_), .Y(n206) );
  XOR3X2_RVT U403 ( .A1(CARRYB_2__8_), .A2(ab_3__8_), .A3(SUMB_2__9_), .Y(
        SUMB_3__8_) );
  NAND2X0_RVT U404 ( .A1(SUMB_2__9_), .A2(CARRYB_2__8_), .Y(n207) );
  NAND2X0_RVT U405 ( .A1(ab_3__8_), .A2(CARRYB_2__8_), .Y(n208) );
  NAND2X0_RVT U406 ( .A1(ab_3__8_), .A2(SUMB_2__9_), .Y(n209) );
  NAND3X0_RVT U407 ( .A1(n209), .A2(n208), .A3(n207), .Y(CARRYB_3__8_) );
  XOR3X2_RVT U408 ( .A1(SUMB_2__10_), .A2(ab_3__9_), .A3(CARRYB_2__9_), .Y(
        SUMB_3__9_) );
  NAND2X0_RVT U409 ( .A1(CARRYB_2__9_), .A2(SUMB_2__10_), .Y(n210) );
  NAND2X0_RVT U410 ( .A1(ab_3__9_), .A2(SUMB_2__10_), .Y(n211) );
  NAND2X0_RVT U411 ( .A1(ab_3__9_), .A2(CARRYB_2__9_), .Y(n212) );
  NAND3X0_RVT U412 ( .A1(n212), .A2(n211), .A3(n210), .Y(CARRYB_3__9_) );
  XOR3X2_RVT U413 ( .A1(n190), .A2(ab_4__21_), .A3(n202), .Y(SUMB_4__21_) );
  NAND2X0_RVT U414 ( .A1(SUMB_3__22_), .A2(n189), .Y(n213) );
  NAND2X0_RVT U415 ( .A1(ab_4__21_), .A2(n189), .Y(n214) );
  NAND2X0_RVT U416 ( .A1(ab_4__21_), .A2(SUMB_3__22_), .Y(n215) );
  NAND3X0_RVT U417 ( .A1(n213), .A2(n215), .A3(n214), .Y(CARRYB_4__21_) );
  AND2X4_RVT U418 ( .A1(n39), .A2(n513), .Y(ab_9__8_) );
  AND2X1_RVT U419 ( .A1(n498), .A2(B[8]), .Y(ab_1__8_) );
  XOR3X2_RVT U420 ( .A1(n173), .A2(ab_5__7_), .A3(n174), .Y(SUMB_5__7_) );
  NAND2X0_RVT U421 ( .A1(CARRYB_4__7_), .A2(SUMB_4__8_), .Y(n216) );
  NAND2X0_RVT U422 ( .A1(ab_5__7_), .A2(CARRYB_4__7_), .Y(n217) );
  NAND2X0_RVT U423 ( .A1(ab_5__7_), .A2(SUMB_4__8_), .Y(n218) );
  NAND3X0_RVT U424 ( .A1(n216), .A2(n218), .A3(n217), .Y(CARRYB_5__7_) );
  AND2X4_RVT U425 ( .A1(n498), .A2(B[4]), .Y(ab_1__4_) );
  AND2X1_RVT U426 ( .A1(n381), .A2(B[9]), .Y(ab_0__9_) );
  NBUFFX2_RVT U427 ( .A(n461), .Y(n220) );
  XOR3X2_RVT U428 ( .A1(CARRYB_25__3_), .A2(ab_26__3_), .A3(SUMB_25__4_), .Y(
        SUMB_26__3_) );
  NAND2X0_RVT U429 ( .A1(SUMB_25__4_), .A2(n169), .Y(n221) );
  NAND2X0_RVT U430 ( .A1(ab_26__3_), .A2(n169), .Y(n222) );
  NAND2X0_RVT U431 ( .A1(ab_26__3_), .A2(SUMB_25__4_), .Y(n223) );
  NBUFFX2_RVT U432 ( .A(n255), .Y(n224) );
  AND2X1_RVT U433 ( .A1(n500), .A2(n255), .Y(ab_3__17_) );
  AND2X1_RVT U434 ( .A1(n503), .A2(n224), .Y(ab_4__17_) );
  NAND3X0_RVT U435 ( .A1(n313), .A2(n314), .A3(n312), .Y(CARRYB_5__12_) );
  XOR2X2_RVT U436 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  XOR3X2_RVT U437 ( .A1(SUMB_5__24_), .A2(ab_6__23_), .A3(CARRYB_5__23_), .Y(
        SUMB_6__23_) );
  NAND2X0_RVT U438 ( .A1(CARRYB_5__23_), .A2(SUMB_5__24_), .Y(n225) );
  NAND2X0_RVT U439 ( .A1(ab_6__23_), .A2(SUMB_5__24_), .Y(n226) );
  NAND2X0_RVT U440 ( .A1(ab_6__23_), .A2(CARRYB_5__23_), .Y(n227) );
  NAND3X0_RVT U441 ( .A1(n227), .A2(n226), .A3(n225), .Y(CARRYB_6__23_) );
  XOR2X1_RVT U442 ( .A1(CARRYB_11__17_), .A2(ab_12__17_), .Y(n228) );
  XOR2X1_RVT U443 ( .A1(n200), .A2(n228), .Y(SUMB_12__17_) );
  AND2X4_RVT U444 ( .A1(n507), .A2(n299), .Y(ab_6__23_) );
  XOR3X2_RVT U445 ( .A1(CARRYB_1__24_), .A2(ab_2__24_), .A3(SUMB_1__25_), .Y(
        n229) );
  XOR2X2_RVT U446 ( .A1(ab_0__24_), .A2(n326), .Y(SUMB_1__23_) );
  NAND3X0_RVT U447 ( .A1(n340), .A2(n341), .A3(n339), .Y(CARRYB_2__20_) );
  AND2X1_RVT U448 ( .A1(B[27]), .A2(n54), .Y(ab_1__27_) );
  AND2X1_RVT U449 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  XOR3X2_RVT U450 ( .A1(SUMB_3__8_), .A2(ab_4__7_), .A3(CARRYB_3__7_), .Y(
        SUMB_4__7_) );
  NAND2X0_RVT U451 ( .A1(CARRYB_3__7_), .A2(SUMB_3__8_), .Y(n230) );
  NAND2X0_RVT U452 ( .A1(ab_4__7_), .A2(SUMB_3__8_), .Y(n231) );
  NAND2X0_RVT U453 ( .A1(ab_4__7_), .A2(CARRYB_3__7_), .Y(n232) );
  NAND3X0_RVT U454 ( .A1(n231), .A2(n232), .A3(n230), .Y(CARRYB_4__7_) );
  AND2X1_RVT U455 ( .A1(n503), .A2(n239), .Y(ab_4__7_) );
  XOR3X2_RVT U456 ( .A1(n144), .A2(ab_6__12_), .A3(SUMB_5__13_), .Y(
        SUMB_6__12_) );
  NAND2X0_RVT U457 ( .A1(SUMB_5__13_), .A2(CARRYB_5__12_), .Y(n233) );
  NAND2X0_RVT U458 ( .A1(ab_6__12_), .A2(CARRYB_5__12_), .Y(n234) );
  NAND2X0_RVT U459 ( .A1(ab_6__12_), .A2(SUMB_5__13_), .Y(n235) );
  NAND3X0_RVT U460 ( .A1(n235), .A2(n234), .A3(n233), .Y(CARRYB_6__12_) );
  NAND2X0_RVT U461 ( .A1(B[22]), .A2(A[0]), .Y(n236) );
  NAND2X0_RVT U462 ( .A1(SUMB_29__1_), .A2(CARRYB_29__0_), .Y(n375) );
  XOR3X2_RVT U463 ( .A1(CARRYB_2__7_), .A2(ab_3__7_), .A3(SUMB_2__8_), .Y(
        SUMB_3__7_) );
  XOR3X2_RVT U464 ( .A1(CARRYB_1__23_), .A2(ab_2__23_), .A3(SUMB_1__24_), .Y(
        SUMB_2__23_) );
  XOR2X1_RVT U465 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  INVX0_RVT U466 ( .A(n495), .Y(n237) );
  IBUFFX8_RVT U467 ( .A(n237), .Y(n238) );
  AND2X1_RVT U468 ( .A1(n248), .A2(B[29]), .Y(ab_2__29_) );
  NBUFFX2_RVT U469 ( .A(n161), .Y(n239) );
  NBUFFX2_RVT U470 ( .A(SUMB_15__14_), .Y(n240) );
  DELLN3X2_RVT U471 ( .A(B[10]), .Y(n455) );
  NAND3X0_RVT U472 ( .A1(n309), .A2(n310), .A3(n311), .Y(n241) );
  NAND3X0_RVT U473 ( .A1(n309), .A2(n310), .A3(n311), .Y(CARRYB_4__15_) );
  NAND3X2_RVT U474 ( .A1(n324), .A2(n323), .A3(n322), .Y(n256) );
  NAND3X2_RVT U475 ( .A1(n305), .A2(n303), .A3(n304), .Y(n247) );
  AND2X1_RVT U476 ( .A1(n501), .A2(n493), .Y(ab_3__6_) );
  NBUFFX2_RVT U477 ( .A(SUMB_3__18_), .Y(n242) );
  NBUFFX2_RVT U478 ( .A(SUMB_23__5_), .Y(n243) );
  AND2X1_RVT U479 ( .A1(A[4]), .A2(n464), .Y(ab_4__22_) );
  XOR2X1_RVT U480 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  AND2X1_RVT U481 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  XOR3X2_RVT U482 ( .A1(ab_13__15_), .A2(CARRYB_12__15_), .A3(SUMB_12__16_), 
        .Y(n244) );
  XOR3X2_RVT U483 ( .A1(ab_8__19_), .A2(CARRYB_7__19_), .A3(SUMB_7__20_), .Y(
        n245) );
  NAND3X0_RVT U484 ( .A1(n303), .A2(n305), .A3(n304), .Y(n246) );
  NAND3X0_RVT U485 ( .A1(n304), .A2(n305), .A3(n303), .Y(CARRYB_2__17_) );
  AND2X1_RVT U486 ( .A1(n501), .A2(n457), .Y(ab_3__12_) );
  NAND2X0_RVT U487 ( .A1(ab_10__19_), .A2(CARRYB_9__19_), .Y(n431) );
  NBUFFX2_RVT U488 ( .A(n499), .Y(n248) );
  NBUFFX2_RVT U489 ( .A(n499), .Y(n249) );
  XOR2X2_RVT U490 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  NBUFFX2_RVT U491 ( .A(n497), .Y(n498) );
  AND2X4_RVT U492 ( .A1(n459), .A2(n512), .Y(ab_9__14_) );
  NAND3X0_RVT U493 ( .A1(n302), .A2(n301), .A3(n300), .Y(n251) );
  AND2X1_RVT U494 ( .A1(n499), .A2(n148), .Y(ab_2__21_) );
  AND2X1_RVT U495 ( .A1(n500), .A2(n148), .Y(ab_3__21_) );
  AND2X1_RVT U496 ( .A1(ab_1__20_), .A2(n138), .Y(CARRYB_1__20_) );
  NAND2X0_RVT U497 ( .A1(ab_7__20_), .A2(CARRYB_6__20_), .Y(n283) );
  AND2X1_RVT U498 ( .A1(n504), .A2(n460), .Y(ab_5__15_) );
  AND2X1_RVT U499 ( .A1(n248), .A2(n460), .Y(ab_2__15_) );
  AND2X1_RVT U500 ( .A1(n501), .A2(n460), .Y(ab_3__15_) );
  XOR3X2_RVT U501 ( .A1(SUMB_2__12_), .A2(ab_3__11_), .A3(CARRYB_2__11_), .Y(
        SUMB_3__11_) );
  NAND2X0_RVT U502 ( .A1(CARRYB_2__11_), .A2(SUMB_2__12_), .Y(n252) );
  NAND2X0_RVT U503 ( .A1(ab_3__11_), .A2(SUMB_2__12_), .Y(n253) );
  NAND2X0_RVT U504 ( .A1(ab_3__11_), .A2(CARRYB_2__11_), .Y(n254) );
  NAND3X0_RVT U505 ( .A1(n254), .A2(n253), .A3(n252), .Y(CARRYB_3__11_) );
  AND2X4_RVT U506 ( .A1(n458), .A2(n512), .Y(ab_9__13_) );
  AND2X1_RVT U507 ( .A1(n502), .A2(n458), .Y(ab_3__13_) );
  NBUFFX2_RVT U508 ( .A(B[17]), .Y(n255) );
  AND2X1_RVT U509 ( .A1(n501), .A2(n220), .Y(ab_3__18_) );
  AND2X1_RVT U510 ( .A1(n499), .A2(n461), .Y(ab_2__18_) );
  XOR3X2_RVT U511 ( .A1(CARRYB_7__20_), .A2(ab_8__20_), .A3(SUMB_7__21_), .Y(
        SUMB_8__20_) );
  NAND2X0_RVT U512 ( .A1(SUMB_7__21_), .A2(n261), .Y(n257) );
  NAND2X0_RVT U513 ( .A1(ab_8__20_), .A2(n261), .Y(n258) );
  NAND2X0_RVT U514 ( .A1(ab_8__20_), .A2(SUMB_7__21_), .Y(n259) );
  NAND3X0_RVT U515 ( .A1(n356), .A2(n355), .A3(n354), .Y(n260) );
  NAND3X0_RVT U516 ( .A1(n283), .A2(n282), .A3(n281), .Y(n261) );
  AND2X1_RVT U517 ( .A1(n499), .A2(B[25]), .Y(ab_2__25_) );
  XOR3X2_RVT U518 ( .A1(SUMB_8__12_), .A2(ab_9__11_), .A3(CARRYB_8__11_), .Y(
        SUMB_9__11_) );
  NAND2X0_RVT U519 ( .A1(CARRYB_8__11_), .A2(SUMB_8__12_), .Y(n262) );
  NAND2X0_RVT U520 ( .A1(ab_9__11_), .A2(SUMB_8__12_), .Y(n263) );
  NAND2X0_RVT U521 ( .A1(ab_9__11_), .A2(CARRYB_8__11_), .Y(n264) );
  NAND3X0_RVT U522 ( .A1(n264), .A2(n263), .A3(n262), .Y(CARRYB_9__11_) );
  XOR3X2_RVT U523 ( .A1(ab_9__20_), .A2(CARRYB_8__20_), .A3(SUMB_8__21_), .Y(
        n265) );
  XOR2X1_RVT U524 ( .A1(CARRYB_18__11_), .A2(ab_19__11_), .Y(n266) );
  XOR2X1_RVT U525 ( .A1(SUMB_18__12_), .A2(n266), .Y(SUMB_19__11_) );
  XOR2X2_RVT U526 ( .A1(ab_0__25_), .A2(n250), .Y(SUMB_1__24_) );
  XOR3X2_RVT U527 ( .A1(CARRYB_2__23_), .A2(ab_3__23_), .A3(SUMB_2__24_), .Y(
        SUMB_3__23_) );
  NAND2X0_RVT U528 ( .A1(n229), .A2(CARRYB_2__23_), .Y(n267) );
  NAND2X0_RVT U529 ( .A1(ab_3__23_), .A2(CARRYB_2__23_), .Y(n268) );
  NAND2X0_RVT U530 ( .A1(ab_3__23_), .A2(n229), .Y(n269) );
  NAND3X0_RVT U531 ( .A1(n269), .A2(n268), .A3(n267), .Y(CARRYB_3__23_) );
  XOR3X2_RVT U532 ( .A1(CARRYB_3__22_), .A2(ab_4__22_), .A3(SUMB_3__23_), .Y(
        SUMB_4__22_) );
  NAND2X0_RVT U533 ( .A1(CARRYB_3__22_), .A2(SUMB_3__23_), .Y(n270) );
  NAND2X0_RVT U534 ( .A1(ab_4__22_), .A2(CARRYB_3__22_), .Y(n271) );
  NAND2X0_RVT U535 ( .A1(ab_4__22_), .A2(SUMB_3__23_), .Y(n272) );
  NAND3X0_RVT U536 ( .A1(n272), .A2(n271), .A3(n270), .Y(CARRYB_4__22_) );
  XOR3X2_RVT U537 ( .A1(SUMB_1__28_), .A2(ab_2__27_), .A3(CARRYB_1__27_), .Y(
        SUMB_2__27_) );
  NAND2X0_RVT U538 ( .A1(CARRYB_1__27_), .A2(SUMB_1__28_), .Y(n273) );
  NAND2X0_RVT U539 ( .A1(ab_2__27_), .A2(SUMB_1__28_), .Y(n274) );
  NAND3X0_RVT U540 ( .A1(n275), .A2(n274), .A3(n273), .Y(CARRYB_2__27_) );
  INVX1_RVT U541 ( .A(n276), .Y(n277) );
  XOR3X2_RVT U542 ( .A1(CARRYB_10__16_), .A2(ab_11__16_), .A3(SUMB_10__17_), 
        .Y(SUMB_11__16_) );
  NAND2X0_RVT U543 ( .A1(SUMB_10__17_), .A2(CARRYB_10__16_), .Y(n278) );
  NAND2X0_RVT U544 ( .A1(ab_11__16_), .A2(CARRYB_10__16_), .Y(n279) );
  NAND2X0_RVT U545 ( .A1(ab_11__16_), .A2(SUMB_10__17_), .Y(n280) );
  NAND3X0_RVT U546 ( .A1(n280), .A2(n279), .A3(n278), .Y(CARRYB_11__16_) );
  XOR3X2_RVT U547 ( .A1(CARRYB_6__20_), .A2(ab_7__20_), .A3(SUMB_6__21_), .Y(
        SUMB_7__20_) );
  NAND2X0_RVT U548 ( .A1(CARRYB_6__20_), .A2(SUMB_6__21_), .Y(n281) );
  NAND2X0_RVT U549 ( .A1(ab_7__20_), .A2(SUMB_6__21_), .Y(n282) );
  NAND3X0_RVT U550 ( .A1(n283), .A2(n282), .A3(n281), .Y(CARRYB_7__20_) );
  NAND2X0_RVT U551 ( .A1(ab_26__2_), .A2(CARRYB_25__2_), .Y(n402) );
  AND2X1_RVT U552 ( .A1(n499), .A2(n463), .Y(ab_2__20_) );
  AND2X1_RVT U553 ( .A1(n504), .A2(n462), .Y(ab_5__19_) );
  AND2X4_RVT U554 ( .A1(n456), .A2(n512), .Y(ab_9__11_) );
  NAND2X0_RVT U555 ( .A1(B[26]), .A2(n381), .Y(n284) );
  XOR3X2_RVT U556 ( .A1(CARRYB_7__11_), .A2(ab_8__11_), .A3(SUMB_7__12_), .Y(
        SUMB_8__11_) );
  NAND2X0_RVT U557 ( .A1(CARRYB_7__11_), .A2(SUMB_7__12_), .Y(n285) );
  NAND2X0_RVT U558 ( .A1(ab_8__11_), .A2(SUMB_7__12_), .Y(n286) );
  NAND2X0_RVT U559 ( .A1(ab_8__11_), .A2(CARRYB_7__11_), .Y(n287) );
  AND2X1_RVT U560 ( .A1(n509), .A2(n464), .Y(ab_7__22_) );
  AND2X1_RVT U561 ( .A1(n499), .A2(n464), .Y(ab_2__22_) );
  AND2X1_RVT U562 ( .A1(n249), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U563 ( .A1(n501), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U564 ( .A1(B[26]), .A2(n325), .Y(n288) );
  XOR3X2_RVT U565 ( .A1(CARRYB_15__13_), .A2(ab_16__13_), .A3(SUMB_15__14_), 
        .Y(SUMB_16__13_) );
  NAND2X0_RVT U566 ( .A1(CARRYB_15__13_), .A2(n240), .Y(n289) );
  NAND2X0_RVT U567 ( .A1(ab_16__13_), .A2(n240), .Y(n290) );
  NAND2X0_RVT U568 ( .A1(ab_16__13_), .A2(CARRYB_15__13_), .Y(n291) );
  NAND3X0_RVT U569 ( .A1(n291), .A2(n290), .A3(n289), .Y(CARRYB_16__13_) );
  NBUFFX2_RVT U570 ( .A(B[15]), .Y(n460) );
  AND2X1_RVT U571 ( .A1(n504), .A2(n457), .Y(ab_5__12_) );
  NAND2X0_RVT U572 ( .A1(ab_5__12_), .A2(CARRYB_4__12_), .Y(n314) );
  XOR3X2_RVT U573 ( .A1(n251), .A2(ab_7__13_), .A3(SUMB_6__14_), .Y(
        SUMB_7__13_) );
  NAND2X0_RVT U574 ( .A1(n251), .A2(SUMB_6__14_), .Y(n292) );
  NAND2X0_RVT U575 ( .A1(ab_7__13_), .A2(SUMB_6__14_), .Y(n293) );
  NAND2X0_RVT U576 ( .A1(ab_7__13_), .A2(n251), .Y(n294) );
  XOR3X2_RVT U577 ( .A1(CARRYB_1__18_), .A2(ab_2__18_), .A3(SUMB_1__19_), .Y(
        SUMB_2__18_) );
  NAND2X0_RVT U578 ( .A1(ab_2__18_), .A2(SUMB_1__19_), .Y(n295) );
  NAND2X0_RVT U579 ( .A1(CARRYB_1__18_), .A2(SUMB_1__19_), .Y(n296) );
  NAND2X0_RVT U580 ( .A1(CARRYB_1__18_), .A2(ab_2__18_), .Y(n297) );
  NAND3X0_RVT U581 ( .A1(n296), .A2(n297), .A3(n295), .Y(CARRYB_2__18_) );
  IBUFFX2_RVT U582 ( .A(B[23]), .Y(n298) );
  INVX1_RVT U583 ( .A(n298), .Y(n299) );
  AND2X1_RVT U584 ( .A1(n505), .A2(n299), .Y(ab_5__23_) );
  XOR3X2_RVT U585 ( .A1(CARRYB_5__13_), .A2(ab_6__13_), .A3(SUMB_5__14_), .Y(
        SUMB_6__13_) );
  NAND2X0_RVT U586 ( .A1(SUMB_5__14_), .A2(CARRYB_5__13_), .Y(n300) );
  NAND2X0_RVT U587 ( .A1(ab_6__13_), .A2(SUMB_5__14_), .Y(n301) );
  NAND2X0_RVT U588 ( .A1(ab_6__13_), .A2(CARRYB_5__13_), .Y(n302) );
  XOR3X2_RVT U589 ( .A1(CARRYB_1__17_), .A2(ab_2__17_), .A3(SUMB_1__18_), .Y(
        SUMB_2__17_) );
  NAND2X0_RVT U590 ( .A1(CARRYB_1__17_), .A2(SUMB_1__18_), .Y(n303) );
  NAND2X0_RVT U591 ( .A1(ab_2__17_), .A2(SUMB_1__18_), .Y(n304) );
  NAND2X0_RVT U592 ( .A1(ab_2__17_), .A2(CARRYB_1__17_), .Y(n305) );
  XOR3X2_RVT U593 ( .A1(ab_2__15_), .A2(CARRYB_1__15_), .A3(SUMB_1__16_), .Y(
        SUMB_2__15_) );
  NAND2X0_RVT U594 ( .A1(ab_2__15_), .A2(SUMB_1__16_), .Y(n306) );
  NAND2X0_RVT U595 ( .A1(CARRYB_1__15_), .A2(ab_2__15_), .Y(n307) );
  NAND2X0_RVT U596 ( .A1(CARRYB_1__15_), .A2(SUMB_1__16_), .Y(n308) );
  XOR2X2_RVT U597 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(SUMB_1__16_) );
  XOR2X2_RVT U598 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR3X2_RVT U599 ( .A1(SUMB_3__16_), .A2(ab_4__15_), .A3(n256), .Y(
        SUMB_4__15_) );
  NAND2X0_RVT U600 ( .A1(SUMB_3__16_), .A2(CARRYB_3__15_), .Y(n309) );
  NAND2X0_RVT U601 ( .A1(ab_4__15_), .A2(SUMB_3__16_), .Y(n310) );
  NAND2X0_RVT U602 ( .A1(ab_4__15_), .A2(n10), .Y(n311) );
  AND2X1_RVT U603 ( .A1(n325), .A2(n461), .Y(ab_0__18_) );
  XOR3X2_RVT U604 ( .A1(CARRYB_4__12_), .A2(ab_5__12_), .A3(SUMB_4__13_), .Y(
        SUMB_5__12_) );
  NAND2X0_RVT U605 ( .A1(CARRYB_4__12_), .A2(SUMB_4__13_), .Y(n312) );
  NAND2X0_RVT U606 ( .A1(ab_5__12_), .A2(SUMB_4__13_), .Y(n313) );
  NBUFFX2_RVT U607 ( .A(SUMB_5__19_), .Y(n315) );
  XOR3X2_RVT U608 ( .A1(n80), .A2(ab_4__17_), .A3(n242), .Y(SUMB_4__17_) );
  NAND2X0_RVT U609 ( .A1(SUMB_3__18_), .A2(CARRYB_3__17_), .Y(n316) );
  NAND2X0_RVT U610 ( .A1(ab_4__17_), .A2(SUMB_3__18_), .Y(n317) );
  NAND2X0_RVT U611 ( .A1(ab_4__17_), .A2(CARRYB_3__17_), .Y(n318) );
  NAND3X0_RVT U612 ( .A1(n316), .A2(n317), .A3(n318), .Y(CARRYB_4__17_) );
  AND2X1_RVT U613 ( .A1(B[26]), .A2(n249), .Y(ab_2__26_) );
  XOR3X2_RVT U614 ( .A1(CARRYB_6__11_), .A2(ab_7__11_), .A3(SUMB_6__12_), .Y(
        SUMB_7__11_) );
  NAND2X0_RVT U615 ( .A1(CARRYB_6__11_), .A2(SUMB_6__12_), .Y(n319) );
  NAND2X0_RVT U616 ( .A1(ab_7__11_), .A2(SUMB_6__12_), .Y(n320) );
  NAND2X0_RVT U617 ( .A1(ab_7__11_), .A2(CARRYB_6__11_), .Y(n321) );
  XOR3X2_RVT U618 ( .A1(n160), .A2(ab_3__15_), .A3(SUMB_2__16_), .Y(
        SUMB_3__15_) );
  NAND2X0_RVT U619 ( .A1(n159), .A2(SUMB_2__16_), .Y(n322) );
  NAND2X0_RVT U620 ( .A1(ab_3__15_), .A2(SUMB_2__16_), .Y(n323) );
  NAND2X0_RVT U621 ( .A1(ab_3__15_), .A2(n159), .Y(n324) );
  NAND3X0_RVT U622 ( .A1(n323), .A2(n324), .A3(n322), .Y(CARRYB_3__15_) );
  NBUFFX2_RVT U623 ( .A(A[0]), .Y(n325) );
  AND2X1_RVT U624 ( .A1(n499), .A2(B[23]), .Y(ab_2__23_) );
  XOR3X2_RVT U625 ( .A1(n241), .A2(ab_5__15_), .A3(SUMB_4__16_), .Y(
        SUMB_5__15_) );
  AND2X4_RVT U626 ( .A1(n457), .A2(n512), .Y(ab_9__12_) );
  AND2X1_RVT U627 ( .A1(B[23]), .A2(A[1]), .Y(n326) );
  AND2X1_RVT U628 ( .A1(n381), .A2(B[12]), .Y(ab_0__12_) );
  XOR3X2_RVT U629 ( .A1(SUMB_2__18_), .A2(ab_3__17_), .A3(n247), .Y(
        SUMB_3__17_) );
  NAND2X0_RVT U630 ( .A1(SUMB_2__18_), .A2(CARRYB_2__17_), .Y(n328) );
  NAND2X0_RVT U631 ( .A1(ab_3__17_), .A2(SUMB_2__18_), .Y(n329) );
  NAND2X0_RVT U632 ( .A1(ab_3__17_), .A2(n246), .Y(n330) );
  NAND3X0_RVT U633 ( .A1(n328), .A2(n329), .A3(n330), .Y(CARRYB_3__17_) );
  IBUFFX2_RVT U634 ( .A(B[26]), .Y(n331) );
  XOR3X2_RVT U635 ( .A1(CARRYB_4__11_), .A2(ab_5__11_), .A3(SUMB_4__12_), .Y(
        SUMB_5__11_) );
  NAND2X0_RVT U636 ( .A1(CARRYB_4__11_), .A2(SUMB_4__12_), .Y(n333) );
  NAND2X0_RVT U637 ( .A1(ab_5__11_), .A2(SUMB_4__12_), .Y(n334) );
  NAND2X0_RVT U638 ( .A1(ab_5__11_), .A2(CARRYB_4__11_), .Y(n335) );
  NAND3X0_RVT U639 ( .A1(n335), .A2(n334), .A3(n333), .Y(CARRYB_5__11_) );
  XOR3X2_RVT U640 ( .A1(SUMB_2__14_), .A2(ab_3__13_), .A3(CARRYB_2__13_), .Y(
        SUMB_3__13_) );
  NAND2X0_RVT U641 ( .A1(CARRYB_2__13_), .A2(SUMB_2__14_), .Y(n336) );
  NAND2X0_RVT U642 ( .A1(ab_3__13_), .A2(SUMB_2__14_), .Y(n337) );
  NAND2X0_RVT U643 ( .A1(ab_3__13_), .A2(CARRYB_2__13_), .Y(n338) );
  NAND3X0_RVT U644 ( .A1(n338), .A2(n337), .A3(n336), .Y(CARRYB_3__13_) );
  XOR3X2_RVT U645 ( .A1(CARRYB_1__20_), .A2(ab_2__20_), .A3(SUMB_1__21_), .Y(
        SUMB_2__20_) );
  NAND2X0_RVT U646 ( .A1(n7), .A2(SUMB_1__21_), .Y(n339) );
  NAND2X0_RVT U647 ( .A1(ab_2__20_), .A2(SUMB_1__21_), .Y(n340) );
  NAND2X0_RVT U648 ( .A1(n7), .A2(ab_2__20_), .Y(n341) );
  INVX0_RVT U649 ( .A(n382), .Y(n383) );
  NAND2X0_RVT U650 ( .A1(ab_24__4_), .A2(CARRYB_23__4_), .Y(n356) );
  XOR3X2_RVT U651 ( .A1(CARRYB_30__0_), .A2(n342), .A3(n343), .Y(PRODUCT_31_)
         );
  NAND2X0_RVT U652 ( .A1(A[31]), .A2(n481), .Y(n342) );
  XOR3X2_RVT U653 ( .A1(SUMB_10__20_), .A2(ab_11__19_), .A3(CARRYB_10__19_), 
        .Y(n344) );
  XOR3X2_RVT U654 ( .A1(CARRYB_2__21_), .A2(ab_3__21_), .A3(n131), .Y(
        SUMB_3__21_) );
  NAND2X0_RVT U655 ( .A1(CARRYB_2__21_), .A2(SUMB_2__22_), .Y(n345) );
  NAND2X0_RVT U656 ( .A1(ab_3__21_), .A2(SUMB_2__22_), .Y(n346) );
  NAND2X0_RVT U657 ( .A1(ab_3__21_), .A2(CARRYB_2__21_), .Y(n347) );
  NAND2X0_RVT U658 ( .A1(n498), .A2(B[25]), .Y(n348) );
  NAND2X0_RVT U659 ( .A1(A[30]), .A2(n483), .Y(n349) );
  AND3X1_RVT U660 ( .A1(n388), .A2(n389), .A3(n387), .Y(n350) );
  AND2X1_RVT U661 ( .A1(n507), .A2(n464), .Y(ab_6__22_) );
  XOR3X2_RVT U662 ( .A1(CARRYB_13__14_), .A2(ab_14__14_), .A3(SUMB_13__15_), 
        .Y(SUMB_14__14_) );
  NAND2X0_RVT U663 ( .A1(n244), .A2(CARRYB_13__14_), .Y(n351) );
  NAND2X0_RVT U664 ( .A1(ab_14__14_), .A2(CARRYB_13__14_), .Y(n352) );
  NAND2X0_RVT U665 ( .A1(ab_14__14_), .A2(n244), .Y(n353) );
  NAND3X0_RVT U666 ( .A1(n353), .A2(n352), .A3(n351), .Y(CARRYB_14__14_) );
  NAND2X0_RVT U667 ( .A1(ab_15__14_), .A2(CARRYB_14__14_), .Y(n421) );
  XOR3X2_RVT U668 ( .A1(CARRYB_23__4_), .A2(ab_24__4_), .A3(n243), .Y(
        SUMB_24__4_) );
  NAND2X0_RVT U669 ( .A1(CARRYB_23__4_), .A2(SUMB_23__5_), .Y(n354) );
  NAND2X0_RVT U670 ( .A1(ab_24__4_), .A2(SUMB_23__5_), .Y(n355) );
  NAND3X0_RVT U671 ( .A1(n355), .A2(n356), .A3(n354), .Y(CARRYB_24__4_) );
  XOR3X2_RVT U672 ( .A1(CARRYB_9__18_), .A2(ab_10__18_), .A3(SUMB_9__19_), .Y(
        SUMB_10__18_) );
  NAND2X0_RVT U673 ( .A1(SUMB_9__19_), .A2(n9), .Y(n357) );
  NAND2X0_RVT U674 ( .A1(ab_10__18_), .A2(n9), .Y(n358) );
  NAND2X0_RVT U675 ( .A1(ab_10__18_), .A2(SUMB_9__19_), .Y(n359) );
  XOR3X2_RVT U676 ( .A1(CARRYB_8__18_), .A2(ab_9__18_), .A3(n245), .Y(
        SUMB_9__18_) );
  NAND2X0_RVT U677 ( .A1(n245), .A2(CARRYB_8__18_), .Y(n360) );
  NAND2X0_RVT U678 ( .A1(ab_9__18_), .A2(CARRYB_8__18_), .Y(n361) );
  NAND2X0_RVT U679 ( .A1(ab_9__18_), .A2(SUMB_8__19_), .Y(n362) );
  XOR3X2_RVT U680 ( .A1(CARRYB_5__18_), .A2(ab_6__18_), .A3(n315), .Y(
        SUMB_6__18_) );
  NAND2X0_RVT U681 ( .A1(SUMB_5__19_), .A2(CARRYB_5__18_), .Y(n363) );
  NAND2X0_RVT U682 ( .A1(ab_6__18_), .A2(CARRYB_5__18_), .Y(n364) );
  NAND2X0_RVT U683 ( .A1(ab_6__18_), .A2(SUMB_5__19_), .Y(n365) );
  XOR3X2_RVT U684 ( .A1(CARRYB_1__19_), .A2(ab_2__19_), .A3(SUMB_1__20_), .Y(
        SUMB_2__19_) );
  NAND2X0_RVT U685 ( .A1(ab_2__19_), .A2(SUMB_1__20_), .Y(n366) );
  NAND2X0_RVT U686 ( .A1(n14), .A2(SUMB_1__20_), .Y(n367) );
  NAND2X0_RVT U687 ( .A1(ab_2__19_), .A2(n14), .Y(n368) );
  NAND3X0_RVT U688 ( .A1(n366), .A2(n368), .A3(n367), .Y(CARRYB_2__19_) );
  XOR3X2_RVT U689 ( .A1(CARRYB_4__19_), .A2(ab_5__19_), .A3(SUMB_4__20_), .Y(
        SUMB_5__19_) );
  NAND2X0_RVT U690 ( .A1(CARRYB_4__19_), .A2(SUMB_4__20_), .Y(n369) );
  NAND2X0_RVT U691 ( .A1(ab_5__19_), .A2(SUMB_4__20_), .Y(n370) );
  NAND2X0_RVT U692 ( .A1(ab_5__19_), .A2(CARRYB_4__19_), .Y(n371) );
  NAND3X0_RVT U693 ( .A1(n370), .A2(n371), .A3(n369), .Y(CARRYB_5__19_) );
  XOR3X2_RVT U694 ( .A1(CARRYB_10__19_), .A2(ab_11__19_), .A3(SUMB_10__20_), 
        .Y(SUMB_11__19_) );
  NAND2X0_RVT U695 ( .A1(CARRYB_10__19_), .A2(SUMB_10__20_), .Y(n372) );
  NAND2X0_RVT U696 ( .A1(ab_11__19_), .A2(SUMB_10__20_), .Y(n373) );
  NAND2X0_RVT U697 ( .A1(ab_11__19_), .A2(CARRYB_10__19_), .Y(n374) );
  NAND3X0_RVT U698 ( .A1(n374), .A2(n373), .A3(n372), .Y(CARRYB_11__19_) );
  XOR3X2_RVT U699 ( .A1(SUMB_29__1_), .A2(ab_30__0_), .A3(n155), .Y(
        PRODUCT_30_) );
  NAND2X0_RVT U700 ( .A1(ab_30__0_), .A2(CARRYB_29__0_), .Y(n376) );
  NAND2X0_RVT U701 ( .A1(ab_30__0_), .A2(SUMB_29__1_), .Y(n377) );
  NAND3X0_RVT U702 ( .A1(n375), .A2(n376), .A3(n377), .Y(CARRYB_30__0_) );
  AND2X1_RVT U703 ( .A1(B[25]), .A2(n53), .Y(ab_1__25_) );
  AND2X4_RVT U704 ( .A1(n54), .A2(B[30]), .Y(ab_1__30_) );
  AND2X4_RVT U705 ( .A1(n53), .A2(B[2]), .Y(ab_1__2_) );
  XOR3X2_RVT U706 ( .A1(SUMB_5__23_), .A2(ab_6__22_), .A3(CARRYB_5__22_), .Y(
        SUMB_6__22_) );
  NAND2X0_RVT U707 ( .A1(CARRYB_5__22_), .A2(SUMB_5__23_), .Y(n378) );
  NAND2X0_RVT U708 ( .A1(ab_6__22_), .A2(SUMB_5__23_), .Y(n379) );
  NAND2X0_RVT U709 ( .A1(ab_6__22_), .A2(CARRYB_5__22_), .Y(n380) );
  NAND2X0_RVT U710 ( .A1(ab_7__22_), .A2(CARRYB_6__22_), .Y(n437) );
  AND2X1_RVT U711 ( .A1(n499), .A2(B[24]), .Y(ab_2__24_) );
  XOR2X2_RVT U712 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  NBUFFX2_RVT U713 ( .A(A[0]), .Y(n381) );
  AND2X4_RVT U714 ( .A1(n57), .A2(n488), .Y(ab_0__3_) );
  IBUFFX2_RVT U715 ( .A(B[25]), .Y(n382) );
  AND2X4_RVT U716 ( .A1(n277), .A2(n513), .Y(ab_9__20_) );
  AND2X1_RVT U717 ( .A1(n500), .A2(n277), .Y(ab_3__20_) );
  XOR3X2_RVT U718 ( .A1(CARRYB_2__20_), .A2(ab_3__20_), .A3(SUMB_2__21_), .Y(
        SUMB_3__20_) );
  NAND2X0_RVT U719 ( .A1(n3), .A2(n29), .Y(n384) );
  NAND2X0_RVT U720 ( .A1(ab_3__20_), .A2(n3), .Y(n385) );
  NAND2X0_RVT U721 ( .A1(ab_3__20_), .A2(n219), .Y(n386) );
  XOR3X2_RVT U722 ( .A1(CARRYB_28__1_), .A2(ab_29__1_), .A3(SUMB_28__2_), .Y(
        SUMB_29__1_) );
  NAND2X0_RVT U723 ( .A1(SUMB_28__2_), .A2(n110), .Y(n387) );
  NAND2X0_RVT U724 ( .A1(ab_29__1_), .A2(SUMB_28__2_), .Y(n388) );
  NAND2X0_RVT U725 ( .A1(ab_29__1_), .A2(n110), .Y(n389) );
  XOR3X2_RVT U726 ( .A1(ab_12__18_), .A2(CARRYB_11__18_), .A3(n344), .Y(n390)
         );
  XOR3X2_RVT U727 ( .A1(CARRYB_3__24_), .A2(ab_4__24_), .A3(SUMB_3__25_), .Y(
        SUMB_4__24_) );
  NAND2X0_RVT U728 ( .A1(CARRYB_3__24_), .A2(SUMB_3__25_), .Y(n391) );
  NAND2X0_RVT U729 ( .A1(ab_4__24_), .A2(SUMB_3__25_), .Y(n392) );
  NAND2X0_RVT U730 ( .A1(ab_4__24_), .A2(CARRYB_3__24_), .Y(n393) );
  XOR3X2_RVT U731 ( .A1(CARRYB_4__23_), .A2(ab_5__23_), .A3(SUMB_4__24_), .Y(
        SUMB_5__23_) );
  NAND2X0_RVT U732 ( .A1(SUMB_4__24_), .A2(CARRYB_4__23_), .Y(n394) );
  NAND2X0_RVT U733 ( .A1(ab_5__23_), .A2(CARRYB_4__23_), .Y(n395) );
  NAND2X0_RVT U734 ( .A1(ab_5__23_), .A2(SUMB_4__24_), .Y(n396) );
  NAND3X0_RVT U735 ( .A1(n396), .A2(n395), .A3(n394), .Y(CARRYB_5__23_) );
  XOR3X2_RVT U736 ( .A1(SUMB_1__27_), .A2(ab_2__26_), .A3(CARRYB_1__26_), .Y(
        SUMB_2__26_) );
  NAND2X0_RVT U737 ( .A1(CARRYB_1__26_), .A2(SUMB_1__27_), .Y(n397) );
  NAND2X0_RVT U738 ( .A1(ab_2__26_), .A2(SUMB_1__27_), .Y(n398) );
  NAND2X0_RVT U739 ( .A1(ab_2__26_), .A2(CARRYB_1__26_), .Y(n399) );
  XOR3X2_RVT U740 ( .A1(CARRYB_25__2_), .A2(ab_26__2_), .A3(SUMB_25__3_), .Y(
        SUMB_26__2_) );
  NAND2X0_RVT U741 ( .A1(CARRYB_25__2_), .A2(SUMB_25__3_), .Y(n400) );
  NAND2X0_RVT U742 ( .A1(ab_26__2_), .A2(SUMB_25__3_), .Y(n401) );
  AND2X4_RVT U743 ( .A1(A[4]), .A2(B[24]), .Y(ab_4__24_) );
  NAND2X0_RVT U744 ( .A1(ab_27__2_), .A2(CARRYB_26__2_), .Y(n434) );
  XOR3X2_RVT U745 ( .A1(CARRYB_24__4_), .A2(ab_25__4_), .A3(SUMB_24__5_), .Y(
        SUMB_25__4_) );
  NAND2X0_RVT U746 ( .A1(SUMB_24__5_), .A2(CARRYB_24__4_), .Y(n403) );
  NAND2X0_RVT U747 ( .A1(ab_25__4_), .A2(SUMB_24__5_), .Y(n404) );
  NAND2X0_RVT U748 ( .A1(ab_25__4_), .A2(n260), .Y(n405) );
  NAND2X0_RVT U749 ( .A1(ab_26__4_), .A2(CARRYB_25__4_), .Y(n452) );
  NAND2X0_RVT U750 ( .A1(ab_27__3_), .A2(CARRYB_26__3_), .Y(n428) );
  NAND2X0_RVT U751 ( .A1(ab_10__20_), .A2(CARRYB_9__20_), .Y(n425) );
  NAND2X0_RVT U752 ( .A1(ab_23__7_), .A2(CARRYB_22__7_), .Y(n412) );
  NAND2X0_RVT U753 ( .A1(ab_19__11_), .A2(CARRYB_18__11_), .Y(n409) );
  NAND2X0_RVT U754 ( .A1(CARRYB_18__11_), .A2(SUMB_18__12_), .Y(n407) );
  NAND2X0_RVT U755 ( .A1(ab_19__11_), .A2(SUMB_18__12_), .Y(n408) );
  NAND3X0_RVT U756 ( .A1(n409), .A2(n408), .A3(n407), .Y(CARRYB_19__11_) );
  NAND2X0_RVT U757 ( .A1(CARRYB_22__7_), .A2(SUMB_22__8_), .Y(n410) );
  NAND2X0_RVT U758 ( .A1(ab_23__7_), .A2(SUMB_22__8_), .Y(n411) );
  NAND3X0_RVT U759 ( .A1(n412), .A2(n411), .A3(n410), .Y(CARRYB_23__7_) );
  XOR3X2_RVT U760 ( .A1(CARRYB_12__17_), .A2(ab_13__17_), .A3(SUMB_12__18_), 
        .Y(SUMB_13__17_) );
  NAND2X0_RVT U761 ( .A1(CARRYB_12__17_), .A2(n390), .Y(n413) );
  NAND2X0_RVT U762 ( .A1(ab_13__17_), .A2(n390), .Y(n414) );
  NAND2X0_RVT U763 ( .A1(ab_13__17_), .A2(CARRYB_12__17_), .Y(n415) );
  NAND3X0_RVT U764 ( .A1(n415), .A2(n414), .A3(n413), .Y(CARRYB_13__17_) );
  NAND2X0_RVT U765 ( .A1(CARRYB_11__17_), .A2(SUMB_11__18_), .Y(n416) );
  NAND2X0_RVT U766 ( .A1(ab_12__17_), .A2(n200), .Y(n417) );
  NAND2X0_RVT U767 ( .A1(ab_12__17_), .A2(CARRYB_11__17_), .Y(n418) );
  XOR3X2_RVT U768 ( .A1(CARRYB_14__14_), .A2(ab_15__14_), .A3(SUMB_14__15_), 
        .Y(SUMB_15__14_) );
  NAND2X0_RVT U769 ( .A1(CARRYB_14__14_), .A2(SUMB_14__15_), .Y(n419) );
  NAND2X0_RVT U770 ( .A1(ab_15__14_), .A2(SUMB_14__15_), .Y(n420) );
  NAND2X0_RVT U771 ( .A1(ab_16__14_), .A2(CARRYB_15__14_), .Y(n443) );
  XOR3X2_RVT U772 ( .A1(CARRYB_26__3_), .A2(ab_27__3_), .A3(SUMB_26__4_), .Y(
        n422) );
  NAND2X0_RVT U773 ( .A1(CARRYB_9__20_), .A2(SUMB_9__21_), .Y(n423) );
  NAND2X0_RVT U774 ( .A1(ab_10__20_), .A2(SUMB_9__21_), .Y(n424) );
  NAND3X0_RVT U775 ( .A1(n425), .A2(n424), .A3(n423), .Y(CARRYB_10__20_) );
  NAND2X0_RVT U776 ( .A1(CARRYB_26__3_), .A2(SUMB_26__4_), .Y(n426) );
  NAND2X0_RVT U777 ( .A1(ab_27__3_), .A2(SUMB_26__4_), .Y(n427) );
  XOR3X2_RVT U778 ( .A1(SUMB_9__20_), .A2(ab_10__19_), .A3(CARRYB_9__19_), .Y(
        SUMB_10__19_) );
  NAND2X0_RVT U779 ( .A1(CARRYB_9__19_), .A2(n265), .Y(n429) );
  NAND2X0_RVT U780 ( .A1(ab_10__19_), .A2(n265), .Y(n430) );
  NAND3X0_RVT U781 ( .A1(n431), .A2(n430), .A3(n429), .Y(CARRYB_10__19_) );
  XOR3X2_RVT U782 ( .A1(SUMB_26__3_), .A2(ab_27__2_), .A3(CARRYB_26__2_), .Y(
        SUMB_27__2_) );
  NAND2X0_RVT U783 ( .A1(CARRYB_26__2_), .A2(n203), .Y(n432) );
  NAND2X0_RVT U784 ( .A1(ab_27__2_), .A2(n203), .Y(n433) );
  XOR3X2_RVT U785 ( .A1(CARRYB_6__22_), .A2(ab_7__22_), .A3(SUMB_6__23_), .Y(
        SUMB_7__22_) );
  NAND2X0_RVT U786 ( .A1(CARRYB_6__22_), .A2(SUMB_6__23_), .Y(n435) );
  NAND2X0_RVT U787 ( .A1(ab_7__22_), .A2(SUMB_6__23_), .Y(n436) );
  NAND2X0_RVT U788 ( .A1(ab_28__2_), .A2(n111), .Y(n440) );
  XOR3X2_RVT U789 ( .A1(CARRYB_27__2_), .A2(ab_28__2_), .A3(n422), .Y(
        SUMB_28__2_) );
  NAND2X0_RVT U790 ( .A1(n111), .A2(n422), .Y(n438) );
  NAND2X0_RVT U791 ( .A1(ab_28__2_), .A2(n422), .Y(n439) );
  XOR3X2_RVT U792 ( .A1(SUMB_15__15_), .A2(ab_16__14_), .A3(CARRYB_15__14_), 
        .Y(SUMB_16__14_) );
  NAND2X0_RVT U793 ( .A1(CARRYB_15__14_), .A2(SUMB_15__15_), .Y(n441) );
  NAND2X0_RVT U794 ( .A1(ab_16__14_), .A2(SUMB_15__15_), .Y(n442) );
  NAND3X0_RVT U795 ( .A1(n443), .A2(n442), .A3(n441), .Y(CARRYB_16__14_) );
  NAND2X0_RVT U796 ( .A1(ab_2__28_), .A2(SUMB_1__29_), .Y(n444) );
  NAND2X0_RVT U797 ( .A1(CARRYB_1__28_), .A2(SUMB_1__29_), .Y(n445) );
  NAND2X0_RVT U798 ( .A1(CARRYB_1__28_), .A2(ab_2__28_), .Y(n446) );
  NAND3X0_RVT U799 ( .A1(n446), .A2(n445), .A3(n444), .Y(CARRYB_2__28_) );
  XOR3X2_RVT U800 ( .A1(CARRYB_2__27_), .A2(ab_3__27_), .A3(SUMB_2__28_), .Y(
        SUMB_3__27_) );
  NAND2X0_RVT U801 ( .A1(CARRYB_2__27_), .A2(SUMB_2__28_), .Y(n447) );
  NAND2X0_RVT U802 ( .A1(ab_3__27_), .A2(SUMB_2__28_), .Y(n448) );
  NAND2X0_RVT U803 ( .A1(ab_3__27_), .A2(CARRYB_2__27_), .Y(n449) );
  NAND3X0_RVT U804 ( .A1(n449), .A2(n448), .A3(n447), .Y(CARRYB_3__27_) );
  XOR3X2_RVT U805 ( .A1(CARRYB_25__4_), .A2(ab_26__4_), .A3(SUMB_25__5_), .Y(
        SUMB_26__4_) );
  NAND2X0_RVT U806 ( .A1(CARRYB_25__4_), .A2(SUMB_25__5_), .Y(n450) );
  NAND2X0_RVT U807 ( .A1(ab_26__4_), .A2(SUMB_25__5_), .Y(n451) );
  NAND3X0_RVT U808 ( .A1(n452), .A2(n451), .A3(n450), .Y(CARRYB_26__4_) );
  AND2X4_RVT U809 ( .A1(n249), .A2(B[28]), .Y(ab_2__28_) );
  XOR2X1_RVT U810 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U811 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U812 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  NBUFFX2_RVT U813 ( .A(B[0]), .Y(n481) );
  NBUFFX2_RVT U814 ( .A(B[9]), .Y(n495) );
  NBUFFX2_RVT U815 ( .A(B[8]), .Y(n494) );
  NBUFFX2_RVT U816 ( .A(A[9]), .Y(n513) );
  NBUFFX2_RVT U817 ( .A(A[9]), .Y(n512) );
  NBUFFX2_RVT U818 ( .A(B[4]), .Y(n489) );
  NBUFFX2_RVT U819 ( .A(B[2]), .Y(n485) );
  NBUFFX2_RVT U820 ( .A(A[5]), .Y(n504) );
  NBUFFX2_RVT U821 ( .A(A[4]), .Y(n503) );
  NBUFFX2_RVT U822 ( .A(A[3]), .Y(n501) );
  NBUFFX2_RVT U823 ( .A(A[3]), .Y(n500) );
  NBUFFX2_RVT U824 ( .A(A[6]), .Y(n506) );
  NBUFFX2_RVT U825 ( .A(A[7]), .Y(n508) );
  NBUFFX2_RVT U826 ( .A(A[7]), .Y(n509) );
  NBUFFX2_RVT U827 ( .A(B[5]), .Y(n491) );
  NBUFFX2_RVT U828 ( .A(B[6]), .Y(n493) );
  NBUFFX2_RVT U829 ( .A(A[8]), .Y(n511) );
  NBUFFX2_RVT U830 ( .A(A[8]), .Y(n510) );
  NBUFFX2_RVT U831 ( .A(B[3]), .Y(n487) );
  NBUFFX2_RVT U832 ( .A(B[1]), .Y(n483) );
  NBUFFX2_RVT U833 ( .A(B[5]), .Y(n492) );
  XNOR3X1_RVT U834 ( .A1(n453), .A2(CARRYB_22__8_), .A3(SUMB_22__9_), .Y(
        SUMB_23__8_) );
  NAND2X0_RVT U835 ( .A1(n480), .A2(n39), .Y(n453) );
  NBUFFX2_RVT U836 ( .A(A[0]), .Y(n496) );
  NBUFFX2_RVT U837 ( .A(A[3]), .Y(n502) );
  NBUFFX2_RVT U838 ( .A(B[0]), .Y(n482) );
  NBUFFX2_RVT U839 ( .A(B[4]), .Y(n490) );
  NBUFFX2_RVT U840 ( .A(B[1]), .Y(n484) );
  NBUFFX2_RVT U841 ( .A(A[5]), .Y(n505) );
  NBUFFX2_RVT U842 ( .A(B[2]), .Y(n486) );
  NBUFFX2_RVT U843 ( .A(A[6]), .Y(n507) );
  NBUFFX2_RVT U844 ( .A(B[3]), .Y(n488) );
  XOR2X1_RVT U845 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  AND2X1_RVT U846 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U847 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U848 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U849 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U850 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U851 ( .A1(n115), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U852 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U853 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U854 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U855 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U856 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U857 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U858 ( .A1(n327), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U859 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U860 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U861 ( .A1(ab_1__23_), .A2(n168), .Y(CARRYB_1__23_) );
  AND2X1_RVT U862 ( .A1(ab_1__25_), .A2(n288), .Y(CARRYB_1__25_) );
  AND2X1_RVT U863 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  XOR2X2_RVT U864 ( .A1(ab_1__28_), .A2(n406), .Y(SUMB_1__28_) );
  AND2X1_RVT U865 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  XOR2X2_RVT U866 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  NBUFFX2_RVT U867 ( .A(A[2]), .Y(n499) );
  AND2X1_RVT U868 ( .A1(B[26]), .A2(n54), .Y(ab_1__26_) );
  AND2X1_RVT U869 ( .A1(n53), .A2(B[28]), .Y(ab_1__28_) );
  NBUFFX2_RVT U870 ( .A(B[10]), .Y(n454) );
  NBUFFX2_RVT U871 ( .A(B[11]), .Y(n456) );
  NBUFFX2_RVT U872 ( .A(B[12]), .Y(n457) );
  NBUFFX2_RVT U873 ( .A(B[13]), .Y(n458) );
  NBUFFX2_RVT U874 ( .A(B[14]), .Y(n459) );
  NBUFFX2_RVT U875 ( .A(B[18]), .Y(n461) );
  NBUFFX2_RVT U876 ( .A(B[20]), .Y(n463) );
  NBUFFX2_RVT U877 ( .A(A[10]), .Y(n465) );
  NBUFFX2_RVT U878 ( .A(A[10]), .Y(n466) );
  NBUFFX2_RVT U879 ( .A(A[11]), .Y(n467) );
  NBUFFX2_RVT U880 ( .A(A[11]), .Y(n468) );
  NBUFFX2_RVT U881 ( .A(A[12]), .Y(n469) );
  NBUFFX2_RVT U882 ( .A(A[13]), .Y(n470) );
  NBUFFX2_RVT U883 ( .A(A[14]), .Y(n471) );
  NBUFFX2_RVT U884 ( .A(A[15]), .Y(n472) );
  NBUFFX2_RVT U885 ( .A(A[16]), .Y(n473) );
  NBUFFX2_RVT U886 ( .A(A[17]), .Y(n474) );
  NBUFFX2_RVT U887 ( .A(A[18]), .Y(n475) );
  NBUFFX2_RVT U888 ( .A(A[19]), .Y(n476) );
  NBUFFX2_RVT U889 ( .A(A[20]), .Y(n477) );
  NBUFFX2_RVT U890 ( .A(A[21]), .Y(n478) );
  NBUFFX2_RVT U891 ( .A(A[22]), .Y(n479) );
  NBUFFX2_RVT U892 ( .A(A[23]), .Y(n480) );
  AND2X1_RVT U893 ( .A1(n238), .A2(n513), .Y(ab_9__9_) );
  AND2X1_RVT U894 ( .A1(n239), .A2(n513), .Y(ab_9__7_) );
  AND2X1_RVT U895 ( .A1(n491), .A2(n513), .Y(ab_9__5_) );
  AND2X1_RVT U896 ( .A1(n490), .A2(n513), .Y(ab_9__4_) );
  AND2X1_RVT U897 ( .A1(n488), .A2(n513), .Y(ab_9__3_) );
  AND2X1_RVT U898 ( .A1(n464), .A2(n513), .Y(ab_9__22_) );
  AND2X1_RVT U899 ( .A1(n462), .A2(n512), .Y(ab_9__19_) );
  AND2X1_RVT U900 ( .A1(n460), .A2(n512), .Y(ab_9__15_) );
  AND2X1_RVT U901 ( .A1(n454), .A2(n512), .Y(ab_9__10_) );
  AND2X1_RVT U902 ( .A1(n481), .A2(n512), .Y(ab_9__0_) );
  AND2X1_RVT U903 ( .A1(n511), .A2(n238), .Y(ab_8__9_) );
  AND2X1_RVT U904 ( .A1(n511), .A2(n494), .Y(ab_8__8_) );
  AND2X1_RVT U905 ( .A1(n511), .A2(n239), .Y(ab_8__7_) );
  AND2X1_RVT U906 ( .A1(n511), .A2(n56), .Y(ab_8__6_) );
  AND2X1_RVT U907 ( .A1(n511), .A2(n491), .Y(ab_8__5_) );
  AND2X1_RVT U908 ( .A1(n511), .A2(n489), .Y(ab_8__4_) );
  AND2X1_RVT U909 ( .A1(n511), .A2(n488), .Y(ab_8__3_) );
  AND2X1_RVT U910 ( .A1(n511), .A2(n485), .Y(ab_8__2_) );
  AND2X1_RVT U911 ( .A1(n511), .A2(n299), .Y(ab_8__23_) );
  AND2X1_RVT U912 ( .A1(n511), .A2(n464), .Y(ab_8__22_) );
  AND2X1_RVT U913 ( .A1(n511), .A2(n148), .Y(ab_8__21_) );
  AND2X1_RVT U914 ( .A1(n511), .A2(n277), .Y(ab_8__20_) );
  AND2X1_RVT U915 ( .A1(n510), .A2(n484), .Y(ab_8__1_) );
  AND2X1_RVT U916 ( .A1(n510), .A2(n462), .Y(ab_8__19_) );
  AND2X1_RVT U917 ( .A1(n510), .A2(n224), .Y(ab_8__17_) );
  AND2X1_RVT U918 ( .A1(n510), .A2(n143), .Y(ab_8__16_) );
  AND2X1_RVT U919 ( .A1(n510), .A2(n460), .Y(ab_8__15_) );
  AND2X1_RVT U920 ( .A1(n510), .A2(n459), .Y(ab_8__14_) );
  AND2X1_RVT U921 ( .A1(n510), .A2(n458), .Y(ab_8__13_) );
  AND2X1_RVT U922 ( .A1(n510), .A2(n457), .Y(ab_8__12_) );
  AND2X1_RVT U923 ( .A1(n510), .A2(n456), .Y(ab_8__11_) );
  AND2X1_RVT U924 ( .A1(n510), .A2(n454), .Y(ab_8__10_) );
  AND2X1_RVT U925 ( .A1(n510), .A2(n481), .Y(ab_8__0_) );
  AND2X1_RVT U926 ( .A1(n509), .A2(n238), .Y(ab_7__9_) );
  AND2X1_RVT U927 ( .A1(n509), .A2(n494), .Y(ab_7__8_) );
  AND2X1_RVT U928 ( .A1(n509), .A2(n239), .Y(ab_7__7_) );
  AND2X1_RVT U929 ( .A1(n509), .A2(n56), .Y(ab_7__6_) );
  AND2X1_RVT U930 ( .A1(n509), .A2(n491), .Y(ab_7__5_) );
  AND2X1_RVT U931 ( .A1(n509), .A2(n489), .Y(ab_7__4_) );
  AND2X1_RVT U932 ( .A1(n509), .A2(n488), .Y(ab_7__3_) );
  AND2X1_RVT U933 ( .A1(n509), .A2(n485), .Y(ab_7__2_) );
  AND2X1_RVT U934 ( .A1(n509), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U935 ( .A1(n509), .A2(n299), .Y(ab_7__23_) );
  AND2X1_RVT U936 ( .A1(n509), .A2(n148), .Y(ab_7__21_) );
  AND2X1_RVT U937 ( .A1(n509), .A2(n277), .Y(ab_7__20_) );
  AND2X1_RVT U938 ( .A1(n508), .A2(n484), .Y(ab_7__1_) );
  AND2X1_RVT U939 ( .A1(n508), .A2(n224), .Y(ab_7__17_) );
  AND2X1_RVT U940 ( .A1(n508), .A2(n143), .Y(ab_7__16_) );
  AND2X1_RVT U941 ( .A1(n508), .A2(n460), .Y(ab_7__15_) );
  AND2X1_RVT U942 ( .A1(n508), .A2(n459), .Y(ab_7__14_) );
  AND2X1_RVT U943 ( .A1(n508), .A2(n458), .Y(ab_7__13_) );
  AND2X1_RVT U944 ( .A1(n508), .A2(n457), .Y(ab_7__12_) );
  AND2X1_RVT U945 ( .A1(n508), .A2(n456), .Y(ab_7__11_) );
  AND2X1_RVT U946 ( .A1(n508), .A2(n454), .Y(ab_7__10_) );
  AND2X1_RVT U947 ( .A1(n508), .A2(n481), .Y(ab_7__0_) );
  AND2X1_RVT U948 ( .A1(n507), .A2(n238), .Y(ab_6__9_) );
  AND2X1_RVT U949 ( .A1(n507), .A2(n494), .Y(ab_6__8_) );
  AND2X1_RVT U950 ( .A1(n507), .A2(n239), .Y(ab_6__7_) );
  AND2X1_RVT U951 ( .A1(n507), .A2(n56), .Y(ab_6__6_) );
  AND2X1_RVT U952 ( .A1(n507), .A2(n491), .Y(ab_6__5_) );
  AND2X1_RVT U953 ( .A1(n507), .A2(n490), .Y(ab_6__4_) );
  AND2X1_RVT U954 ( .A1(n507), .A2(n488), .Y(ab_6__3_) );
  AND2X1_RVT U955 ( .A1(n507), .A2(n485), .Y(ab_6__2_) );
  AND2X1_RVT U956 ( .A1(n507), .A2(n383), .Y(ab_6__25_) );
  AND2X1_RVT U957 ( .A1(n507), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U958 ( .A1(n506), .A2(n277), .Y(ab_6__20_) );
  AND2X1_RVT U959 ( .A1(n507), .A2(n484), .Y(ab_6__1_) );
  AND2X1_RVT U960 ( .A1(n506), .A2(n462), .Y(ab_6__19_) );
  AND2X1_RVT U961 ( .A1(n506), .A2(n220), .Y(ab_6__18_) );
  AND2X1_RVT U962 ( .A1(n506), .A2(n224), .Y(ab_6__17_) );
  AND2X1_RVT U963 ( .A1(n506), .A2(n143), .Y(ab_6__16_) );
  AND2X1_RVT U964 ( .A1(n507), .A2(n460), .Y(ab_6__15_) );
  AND2X1_RVT U965 ( .A1(n507), .A2(n459), .Y(ab_6__14_) );
  AND2X1_RVT U966 ( .A1(n507), .A2(n458), .Y(ab_6__13_) );
  AND2X1_RVT U967 ( .A1(n507), .A2(n456), .Y(ab_6__11_) );
  AND2X1_RVT U968 ( .A1(n507), .A2(n454), .Y(ab_6__10_) );
  AND2X1_RVT U969 ( .A1(n507), .A2(n481), .Y(ab_6__0_) );
  AND2X1_RVT U970 ( .A1(n505), .A2(n494), .Y(ab_5__8_) );
  AND2X1_RVT U971 ( .A1(n505), .A2(n239), .Y(ab_5__7_) );
  AND2X1_RVT U972 ( .A1(n505), .A2(n56), .Y(ab_5__6_) );
  AND2X1_RVT U973 ( .A1(n505), .A2(n491), .Y(ab_5__5_) );
  AND2X1_RVT U974 ( .A1(n505), .A2(n489), .Y(ab_5__4_) );
  AND2X1_RVT U975 ( .A1(n505), .A2(n488), .Y(ab_5__3_) );
  AND2X1_RVT U976 ( .A1(n505), .A2(n485), .Y(ab_5__2_) );
  AND2X1_RVT U977 ( .A1(n504), .A2(n332), .Y(ab_5__26_) );
  AND2X1_RVT U978 ( .A1(n505), .A2(n383), .Y(ab_5__25_) );
  AND2X1_RVT U979 ( .A1(n505), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U980 ( .A1(n505), .A2(n464), .Y(ab_5__22_) );
  AND2X1_RVT U981 ( .A1(n505), .A2(n277), .Y(ab_5__20_) );
  AND2X1_RVT U982 ( .A1(n504), .A2(n484), .Y(ab_5__1_) );
  AND2X1_RVT U983 ( .A1(n504), .A2(n220), .Y(ab_5__18_) );
  AND2X1_RVT U984 ( .A1(n504), .A2(n224), .Y(ab_5__17_) );
  AND2X1_RVT U985 ( .A1(n504), .A2(n143), .Y(ab_5__16_) );
  AND2X1_RVT U986 ( .A1(n504), .A2(n459), .Y(ab_5__14_) );
  AND2X1_RVT U987 ( .A1(n504), .A2(n458), .Y(ab_5__13_) );
  AND2X1_RVT U988 ( .A1(n504), .A2(n456), .Y(ab_5__11_) );
  AND2X1_RVT U989 ( .A1(n504), .A2(n454), .Y(ab_5__10_) );
  AND2X1_RVT U990 ( .A1(n504), .A2(n481), .Y(ab_5__0_) );
  AND2X1_RVT U991 ( .A1(n503), .A2(n238), .Y(ab_4__9_) );
  AND2X1_RVT U992 ( .A1(n503), .A2(n494), .Y(ab_4__8_) );
  AND2X1_RVT U993 ( .A1(A[4]), .A2(n491), .Y(ab_4__5_) );
  AND2X1_RVT U994 ( .A1(A[4]), .A2(n490), .Y(ab_4__4_) );
  AND2X1_RVT U995 ( .A1(A[4]), .A2(n488), .Y(ab_4__3_) );
  AND2X1_RVT U996 ( .A1(A[4]), .A2(n485), .Y(ab_4__2_) );
  AND2X1_RVT U997 ( .A1(A[4]), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U998 ( .A1(A[4]), .A2(n332), .Y(ab_4__26_) );
  AND2X1_RVT U999 ( .A1(A[4]), .A2(n383), .Y(ab_4__25_) );
  AND2X1_RVT U1000 ( .A1(A[4]), .A2(n299), .Y(ab_4__23_) );
  AND2X1_RVT U1001 ( .A1(A[4]), .A2(n148), .Y(ab_4__21_) );
  AND2X1_RVT U1002 ( .A1(A[4]), .A2(n277), .Y(ab_4__20_) );
  AND2X1_RVT U1003 ( .A1(n503), .A2(n484), .Y(ab_4__1_) );
  AND2X1_RVT U1004 ( .A1(n503), .A2(n220), .Y(ab_4__18_) );
  AND2X1_RVT U1005 ( .A1(n503), .A2(n143), .Y(ab_4__16_) );
  AND2X1_RVT U1006 ( .A1(n503), .A2(n460), .Y(ab_4__15_) );
  AND2X1_RVT U1007 ( .A1(n503), .A2(n459), .Y(ab_4__14_) );
  AND2X1_RVT U1008 ( .A1(n503), .A2(n458), .Y(ab_4__13_) );
  AND2X1_RVT U1009 ( .A1(n503), .A2(n457), .Y(ab_4__12_) );
  AND2X1_RVT U1010 ( .A1(n503), .A2(n456), .Y(ab_4__11_) );
  AND2X1_RVT U1011 ( .A1(n503), .A2(n454), .Y(ab_4__10_) );
  AND2X1_RVT U1012 ( .A1(n503), .A2(n481), .Y(ab_4__0_) );
  AND2X1_RVT U1013 ( .A1(n500), .A2(n494), .Y(ab_3__8_) );
  AND2X1_RVT U1014 ( .A1(n502), .A2(n239), .Y(ab_3__7_) );
  AND2X1_RVT U1015 ( .A1(n500), .A2(n491), .Y(ab_3__5_) );
  AND2X1_RVT U1016 ( .A1(n502), .A2(n489), .Y(ab_3__4_) );
  AND2X1_RVT U1017 ( .A1(n500), .A2(n485), .Y(ab_3__2_) );
  AND2X1_RVT U1018 ( .A1(n500), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U1019 ( .A1(n500), .A2(n332), .Y(ab_3__26_) );
  AND2X1_RVT U1020 ( .A1(n502), .A2(n383), .Y(ab_3__25_) );
  AND2X1_RVT U1021 ( .A1(n502), .A2(n464), .Y(ab_3__22_) );
  AND2X1_RVT U1022 ( .A1(n502), .A2(n484), .Y(ab_3__1_) );
  AND2X1_RVT U1023 ( .A1(n502), .A2(n462), .Y(ab_3__19_) );
  AND2X1_RVT U1024 ( .A1(n502), .A2(n143), .Y(ab_3__16_) );
  AND2X1_RVT U1025 ( .A1(n500), .A2(n459), .Y(ab_3__14_) );
  AND2X1_RVT U1026 ( .A1(n500), .A2(n456), .Y(ab_3__11_) );
  AND2X1_RVT U1027 ( .A1(n502), .A2(n454), .Y(ab_3__10_) );
  AND2X1_RVT U1028 ( .A1(A[30]), .A2(n481), .Y(ab_30__0_) );
  AND2X1_RVT U1029 ( .A1(n248), .A2(n495), .Y(ab_2__9_) );
  AND2X1_RVT U1030 ( .A1(n249), .A2(n494), .Y(ab_2__8_) );
  AND2X1_RVT U1031 ( .A1(n248), .A2(n161), .Y(ab_2__7_) );
  AND2X1_RVT U1032 ( .A1(n248), .A2(n493), .Y(ab_2__6_) );
  AND2X1_RVT U1033 ( .A1(n249), .A2(n491), .Y(ab_2__5_) );
  AND2X1_RVT U1034 ( .A1(n248), .A2(n484), .Y(ab_2__1_) );
  AND2X1_RVT U1035 ( .A1(n499), .A2(B[19]), .Y(ab_2__19_) );
  AND2X1_RVT U1036 ( .A1(n499), .A2(n255), .Y(ab_2__17_) );
  AND2X1_RVT U1037 ( .A1(n249), .A2(B[16]), .Y(ab_2__16_) );
  AND2X1_RVT U1038 ( .A1(n249), .A2(n459), .Y(ab_2__14_) );
  AND2X1_RVT U1039 ( .A1(n248), .A2(n458), .Y(ab_2__13_) );
  AND2X1_RVT U1040 ( .A1(n249), .A2(n457), .Y(ab_2__12_) );
  AND2X1_RVT U1041 ( .A1(n248), .A2(n456), .Y(ab_2__11_) );
  AND2X1_RVT U1042 ( .A1(n249), .A2(n454), .Y(ab_2__10_) );
  AND2X1_RVT U1043 ( .A1(n249), .A2(n481), .Y(ab_2__0_) );
  AND2X1_RVT U1044 ( .A1(A[29]), .A2(n484), .Y(ab_29__1_) );
  AND2X1_RVT U1045 ( .A1(A[29]), .A2(n481), .Y(ab_29__0_) );
  AND2X1_RVT U1046 ( .A1(A[28]), .A2(n485), .Y(ab_28__2_) );
  AND2X1_RVT U1047 ( .A1(A[28]), .A2(n484), .Y(ab_28__1_) );
  AND2X1_RVT U1048 ( .A1(A[28]), .A2(n481), .Y(ab_28__0_) );
  AND2X1_RVT U1049 ( .A1(A[27]), .A2(n490), .Y(ab_27__4_) );
  AND2X1_RVT U1050 ( .A1(A[27]), .A2(n488), .Y(ab_27__3_) );
  AND2X1_RVT U1051 ( .A1(A[27]), .A2(n485), .Y(ab_27__2_) );
  AND2X1_RVT U1052 ( .A1(A[27]), .A2(n484), .Y(ab_27__1_) );
  AND2X1_RVT U1053 ( .A1(A[27]), .A2(n481), .Y(ab_27__0_) );
  AND2X1_RVT U1054 ( .A1(A[26]), .A2(n491), .Y(ab_26__5_) );
  AND2X1_RVT U1055 ( .A1(A[26]), .A2(n489), .Y(ab_26__4_) );
  AND2X1_RVT U1056 ( .A1(A[26]), .A2(n488), .Y(ab_26__3_) );
  AND2X1_RVT U1057 ( .A1(A[26]), .A2(n485), .Y(ab_26__2_) );
  AND2X1_RVT U1058 ( .A1(A[26]), .A2(n484), .Y(ab_26__1_) );
  AND2X1_RVT U1059 ( .A1(A[26]), .A2(n482), .Y(ab_26__0_) );
  AND2X1_RVT U1060 ( .A1(A[25]), .A2(n56), .Y(ab_25__6_) );
  AND2X1_RVT U1061 ( .A1(A[25]), .A2(n491), .Y(ab_25__5_) );
  AND2X1_RVT U1062 ( .A1(A[25]), .A2(n490), .Y(ab_25__4_) );
  AND2X1_RVT U1063 ( .A1(A[25]), .A2(n488), .Y(ab_25__3_) );
  AND2X1_RVT U1064 ( .A1(A[25]), .A2(n485), .Y(ab_25__2_) );
  AND2X1_RVT U1065 ( .A1(A[25]), .A2(n483), .Y(ab_25__1_) );
  AND2X1_RVT U1066 ( .A1(A[25]), .A2(n482), .Y(ab_25__0_) );
  AND2X1_RVT U1067 ( .A1(A[24]), .A2(n239), .Y(ab_24__7_) );
  AND2X1_RVT U1068 ( .A1(A[24]), .A2(n56), .Y(ab_24__6_) );
  AND2X1_RVT U1069 ( .A1(A[24]), .A2(n491), .Y(ab_24__5_) );
  AND2X1_RVT U1070 ( .A1(A[24]), .A2(n489), .Y(ab_24__4_) );
  AND2X1_RVT U1071 ( .A1(A[24]), .A2(n488), .Y(ab_24__3_) );
  AND2X1_RVT U1072 ( .A1(A[24]), .A2(n485), .Y(ab_24__2_) );
  AND2X1_RVT U1073 ( .A1(A[24]), .A2(n483), .Y(ab_24__1_) );
  AND2X1_RVT U1074 ( .A1(A[24]), .A2(n482), .Y(ab_24__0_) );
  AND2X1_RVT U1075 ( .A1(n480), .A2(n239), .Y(ab_23__7_) );
  AND2X1_RVT U1076 ( .A1(n480), .A2(n56), .Y(ab_23__6_) );
  AND2X1_RVT U1077 ( .A1(A[23]), .A2(n491), .Y(ab_23__5_) );
  AND2X1_RVT U1078 ( .A1(n480), .A2(n490), .Y(ab_23__4_) );
  AND2X1_RVT U1079 ( .A1(n480), .A2(n487), .Y(ab_23__3_) );
  AND2X1_RVT U1080 ( .A1(n480), .A2(n486), .Y(ab_23__2_) );
  AND2X1_RVT U1081 ( .A1(n480), .A2(n483), .Y(ab_23__1_) );
  AND2X1_RVT U1082 ( .A1(n480), .A2(n482), .Y(ab_23__0_) );
  AND2X1_RVT U1083 ( .A1(n479), .A2(n238), .Y(ab_22__9_) );
  AND2X1_RVT U1084 ( .A1(n479), .A2(n39), .Y(ab_22__8_) );
  AND2X1_RVT U1085 ( .A1(n479), .A2(n239), .Y(ab_22__7_) );
  AND2X1_RVT U1086 ( .A1(A[22]), .A2(n56), .Y(ab_22__6_) );
  AND2X1_RVT U1087 ( .A1(n479), .A2(n491), .Y(ab_22__5_) );
  AND2X1_RVT U1088 ( .A1(n479), .A2(n489), .Y(ab_22__4_) );
  AND2X1_RVT U1089 ( .A1(n479), .A2(n487), .Y(ab_22__3_) );
  AND2X1_RVT U1090 ( .A1(n479), .A2(n486), .Y(ab_22__2_) );
  AND2X1_RVT U1091 ( .A1(n479), .A2(n483), .Y(ab_22__1_) );
  AND2X1_RVT U1092 ( .A1(n479), .A2(n482), .Y(ab_22__0_) );
  AND2X1_RVT U1093 ( .A1(n478), .A2(n238), .Y(ab_21__9_) );
  AND2X1_RVT U1094 ( .A1(n478), .A2(n39), .Y(ab_21__8_) );
  AND2X1_RVT U1095 ( .A1(n478), .A2(n239), .Y(ab_21__7_) );
  AND2X1_RVT U1096 ( .A1(n478), .A2(n56), .Y(ab_21__6_) );
  AND2X1_RVT U1097 ( .A1(n478), .A2(n492), .Y(ab_21__5_) );
  AND2X1_RVT U1098 ( .A1(n478), .A2(n490), .Y(ab_21__4_) );
  AND2X1_RVT U1099 ( .A1(n478), .A2(n487), .Y(ab_21__3_) );
  AND2X1_RVT U1100 ( .A1(n478), .A2(n486), .Y(ab_21__2_) );
  AND2X1_RVT U1101 ( .A1(n478), .A2(n483), .Y(ab_21__1_) );
  AND2X1_RVT U1102 ( .A1(A[21]), .A2(n454), .Y(ab_21__10_) );
  AND2X1_RVT U1103 ( .A1(n478), .A2(n482), .Y(ab_21__0_) );
  AND2X1_RVT U1104 ( .A1(n477), .A2(n238), .Y(ab_20__9_) );
  AND2X1_RVT U1105 ( .A1(n477), .A2(n39), .Y(ab_20__8_) );
  AND2X1_RVT U1106 ( .A1(n477), .A2(n239), .Y(ab_20__7_) );
  AND2X1_RVT U1107 ( .A1(n477), .A2(n56), .Y(ab_20__6_) );
  AND2X1_RVT U1108 ( .A1(n477), .A2(n492), .Y(ab_20__5_) );
  AND2X1_RVT U1109 ( .A1(n477), .A2(n489), .Y(ab_20__4_) );
  AND2X1_RVT U1110 ( .A1(n477), .A2(n487), .Y(ab_20__3_) );
  AND2X1_RVT U1111 ( .A1(n477), .A2(n486), .Y(ab_20__2_) );
  AND2X1_RVT U1112 ( .A1(n477), .A2(n483), .Y(ab_20__1_) );
  AND2X1_RVT U1113 ( .A1(n477), .A2(n24), .Y(ab_20__11_) );
  AND2X1_RVT U1114 ( .A1(n477), .A2(n454), .Y(ab_20__10_) );
  AND2X1_RVT U1115 ( .A1(n477), .A2(n482), .Y(ab_20__0_) );
  AND2X1_RVT U1116 ( .A1(n498), .A2(B[9]), .Y(ab_1__9_) );
  AND2X1_RVT U1117 ( .A1(n498), .A2(n161), .Y(ab_1__7_) );
  AND2X1_RVT U1118 ( .A1(n498), .A2(B[6]), .Y(ab_1__6_) );
  AND2X1_RVT U1119 ( .A1(n497), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U1120 ( .A1(n461), .A2(n497), .Y(ab_1__18_) );
  AND2X1_RVT U1121 ( .A1(n53), .A2(B[17]), .Y(ab_1__17_) );
  AND2X1_RVT U1122 ( .A1(n54), .A2(B[14]), .Y(ab_1__14_) );
  AND2X1_RVT U1123 ( .A1(n54), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U1124 ( .A1(n54), .A2(B[11]), .Y(ab_1__11_) );
  AND2X1_RVT U1125 ( .A1(n476), .A2(n238), .Y(ab_19__9_) );
  AND2X1_RVT U1126 ( .A1(n476), .A2(n39), .Y(ab_19__8_) );
  AND2X1_RVT U1127 ( .A1(n476), .A2(n239), .Y(ab_19__7_) );
  AND2X1_RVT U1128 ( .A1(n476), .A2(n56), .Y(ab_19__6_) );
  AND2X1_RVT U1129 ( .A1(n476), .A2(n492), .Y(ab_19__5_) );
  AND2X1_RVT U1130 ( .A1(n476), .A2(n490), .Y(ab_19__4_) );
  AND2X1_RVT U1131 ( .A1(n476), .A2(n487), .Y(ab_19__3_) );
  AND2X1_RVT U1132 ( .A1(n476), .A2(n486), .Y(ab_19__2_) );
  AND2X1_RVT U1133 ( .A1(n476), .A2(n483), .Y(ab_19__1_) );
  AND2X1_RVT U1134 ( .A1(n476), .A2(n457), .Y(ab_19__12_) );
  AND2X1_RVT U1135 ( .A1(n476), .A2(n24), .Y(ab_19__11_) );
  AND2X1_RVT U1136 ( .A1(n476), .A2(n455), .Y(ab_19__10_) );
  AND2X1_RVT U1137 ( .A1(n476), .A2(n482), .Y(ab_19__0_) );
  AND2X1_RVT U1138 ( .A1(n475), .A2(n238), .Y(ab_18__9_) );
  AND2X1_RVT U1139 ( .A1(n475), .A2(n39), .Y(ab_18__8_) );
  AND2X1_RVT U1140 ( .A1(n475), .A2(n239), .Y(ab_18__7_) );
  AND2X1_RVT U1141 ( .A1(n475), .A2(n56), .Y(ab_18__6_) );
  AND2X1_RVT U1142 ( .A1(n475), .A2(n492), .Y(ab_18__5_) );
  AND2X1_RVT U1143 ( .A1(n475), .A2(n489), .Y(ab_18__4_) );
  AND2X1_RVT U1144 ( .A1(n475), .A2(n487), .Y(ab_18__3_) );
  AND2X1_RVT U1145 ( .A1(n475), .A2(n486), .Y(ab_18__2_) );
  AND2X1_RVT U1146 ( .A1(n475), .A2(n483), .Y(ab_18__1_) );
  AND2X1_RVT U1147 ( .A1(A[18]), .A2(n458), .Y(ab_18__13_) );
  AND2X1_RVT U1148 ( .A1(n475), .A2(n457), .Y(ab_18__12_) );
  AND2X1_RVT U1149 ( .A1(n475), .A2(n24), .Y(ab_18__11_) );
  AND2X1_RVT U1150 ( .A1(n475), .A2(n455), .Y(ab_18__10_) );
  AND2X1_RVT U1151 ( .A1(n475), .A2(n482), .Y(ab_18__0_) );
  AND2X1_RVT U1152 ( .A1(n474), .A2(n238), .Y(ab_17__9_) );
  AND2X1_RVT U1153 ( .A1(n474), .A2(n39), .Y(ab_17__8_) );
  AND2X1_RVT U1154 ( .A1(n474), .A2(n239), .Y(ab_17__7_) );
  AND2X1_RVT U1155 ( .A1(n474), .A2(n56), .Y(ab_17__6_) );
  AND2X1_RVT U1156 ( .A1(n474), .A2(n492), .Y(ab_17__5_) );
  AND2X1_RVT U1157 ( .A1(n474), .A2(n490), .Y(ab_17__4_) );
  AND2X1_RVT U1158 ( .A1(n474), .A2(n487), .Y(ab_17__3_) );
  AND2X1_RVT U1159 ( .A1(n474), .A2(n486), .Y(ab_17__2_) );
  AND2X1_RVT U1160 ( .A1(n474), .A2(n483), .Y(ab_17__1_) );
  AND2X1_RVT U1161 ( .A1(A[17]), .A2(n5), .Y(ab_17__14_) );
  AND2X1_RVT U1162 ( .A1(n474), .A2(n458), .Y(ab_17__13_) );
  AND2X1_RVT U1163 ( .A1(n474), .A2(n457), .Y(ab_17__12_) );
  AND2X1_RVT U1164 ( .A1(n474), .A2(n24), .Y(ab_17__11_) );
  AND2X1_RVT U1165 ( .A1(A[17]), .A2(n455), .Y(ab_17__10_) );
  AND2X1_RVT U1166 ( .A1(n474), .A2(n482), .Y(ab_17__0_) );
  AND2X1_RVT U1167 ( .A1(n473), .A2(n238), .Y(ab_16__9_) );
  AND2X1_RVT U1168 ( .A1(n473), .A2(n39), .Y(ab_16__8_) );
  AND2X1_RVT U1169 ( .A1(n473), .A2(n239), .Y(ab_16__7_) );
  AND2X1_RVT U1170 ( .A1(n473), .A2(n56), .Y(ab_16__6_) );
  AND2X1_RVT U1171 ( .A1(n473), .A2(n492), .Y(ab_16__5_) );
  AND2X1_RVT U1172 ( .A1(n473), .A2(n489), .Y(ab_16__4_) );
  AND2X1_RVT U1173 ( .A1(n473), .A2(n487), .Y(ab_16__3_) );
  AND2X1_RVT U1174 ( .A1(n473), .A2(n486), .Y(ab_16__2_) );
  AND2X1_RVT U1175 ( .A1(n473), .A2(n483), .Y(ab_16__1_) );
  AND2X1_RVT U1176 ( .A1(A[16]), .A2(n460), .Y(ab_16__15_) );
  AND2X1_RVT U1177 ( .A1(n473), .A2(n5), .Y(ab_16__14_) );
  AND2X1_RVT U1178 ( .A1(n473), .A2(n458), .Y(ab_16__13_) );
  AND2X1_RVT U1179 ( .A1(n473), .A2(n457), .Y(ab_16__12_) );
  AND2X1_RVT U1180 ( .A1(A[16]), .A2(n24), .Y(ab_16__11_) );
  AND2X1_RVT U1181 ( .A1(n473), .A2(n455), .Y(ab_16__10_) );
  AND2X1_RVT U1182 ( .A1(n473), .A2(n482), .Y(ab_16__0_) );
  AND2X1_RVT U1183 ( .A1(n472), .A2(n238), .Y(ab_15__9_) );
  AND2X1_RVT U1184 ( .A1(n472), .A2(n39), .Y(ab_15__8_) );
  AND2X1_RVT U1185 ( .A1(n472), .A2(n239), .Y(ab_15__7_) );
  AND2X1_RVT U1186 ( .A1(n472), .A2(n56), .Y(ab_15__6_) );
  AND2X1_RVT U1187 ( .A1(n472), .A2(n492), .Y(ab_15__5_) );
  AND2X1_RVT U1188 ( .A1(n472), .A2(n490), .Y(ab_15__4_) );
  AND2X1_RVT U1189 ( .A1(A[15]), .A2(n487), .Y(ab_15__3_) );
  AND2X1_RVT U1190 ( .A1(n472), .A2(n486), .Y(ab_15__2_) );
  AND2X1_RVT U1191 ( .A1(A[15]), .A2(n483), .Y(ab_15__1_) );
  AND2X1_RVT U1192 ( .A1(n472), .A2(n143), .Y(ab_15__16_) );
  AND2X1_RVT U1193 ( .A1(n472), .A2(n460), .Y(ab_15__15_) );
  AND2X1_RVT U1194 ( .A1(n472), .A2(n5), .Y(ab_15__14_) );
  AND2X1_RVT U1195 ( .A1(n472), .A2(n458), .Y(ab_15__13_) );
  AND2X1_RVT U1196 ( .A1(n472), .A2(n457), .Y(ab_15__12_) );
  AND2X1_RVT U1197 ( .A1(n472), .A2(n24), .Y(ab_15__11_) );
  AND2X1_RVT U1198 ( .A1(n472), .A2(n455), .Y(ab_15__10_) );
  AND2X1_RVT U1199 ( .A1(A[15]), .A2(n482), .Y(ab_15__0_) );
  AND2X1_RVT U1200 ( .A1(n471), .A2(n238), .Y(ab_14__9_) );
  AND2X1_RVT U1201 ( .A1(n471), .A2(n39), .Y(ab_14__8_) );
  AND2X1_RVT U1202 ( .A1(n471), .A2(n239), .Y(ab_14__7_) );
  AND2X1_RVT U1203 ( .A1(n471), .A2(n56), .Y(ab_14__6_) );
  AND2X1_RVT U1204 ( .A1(n471), .A2(n492), .Y(ab_14__5_) );
  AND2X1_RVT U1205 ( .A1(n471), .A2(n489), .Y(ab_14__4_) );
  AND2X1_RVT U1206 ( .A1(n471), .A2(n487), .Y(ab_14__3_) );
  AND2X1_RVT U1207 ( .A1(A[14]), .A2(n486), .Y(ab_14__2_) );
  AND2X1_RVT U1208 ( .A1(n471), .A2(n483), .Y(ab_14__1_) );
  AND2X1_RVT U1209 ( .A1(A[14]), .A2(n224), .Y(ab_14__17_) );
  AND2X1_RVT U1210 ( .A1(n471), .A2(n143), .Y(ab_14__16_) );
  AND2X1_RVT U1211 ( .A1(n471), .A2(n460), .Y(ab_14__15_) );
  AND2X1_RVT U1212 ( .A1(n471), .A2(n5), .Y(ab_14__14_) );
  AND2X1_RVT U1213 ( .A1(A[14]), .A2(n458), .Y(ab_14__13_) );
  AND2X1_RVT U1214 ( .A1(n471), .A2(n457), .Y(ab_14__12_) );
  AND2X1_RVT U1215 ( .A1(n471), .A2(n24), .Y(ab_14__11_) );
  AND2X1_RVT U1216 ( .A1(n471), .A2(n455), .Y(ab_14__10_) );
  AND2X1_RVT U1217 ( .A1(A[14]), .A2(n482), .Y(ab_14__0_) );
  AND2X1_RVT U1218 ( .A1(n470), .A2(n238), .Y(ab_13__9_) );
  AND2X1_RVT U1219 ( .A1(n470), .A2(n39), .Y(ab_13__8_) );
  AND2X1_RVT U1220 ( .A1(n470), .A2(n239), .Y(ab_13__7_) );
  AND2X1_RVT U1221 ( .A1(A[13]), .A2(n56), .Y(ab_13__6_) );
  AND2X1_RVT U1222 ( .A1(n470), .A2(n492), .Y(ab_13__5_) );
  AND2X1_RVT U1223 ( .A1(A[13]), .A2(n490), .Y(ab_13__4_) );
  AND2X1_RVT U1224 ( .A1(n470), .A2(n487), .Y(ab_13__3_) );
  AND2X1_RVT U1225 ( .A1(A[13]), .A2(n486), .Y(ab_13__2_) );
  AND2X1_RVT U1226 ( .A1(n470), .A2(n483), .Y(ab_13__1_) );
  AND2X1_RVT U1227 ( .A1(A[13]), .A2(n220), .Y(ab_13__18_) );
  AND2X1_RVT U1228 ( .A1(n470), .A2(n224), .Y(ab_13__17_) );
  AND2X1_RVT U1229 ( .A1(n470), .A2(n143), .Y(ab_13__16_) );
  AND2X1_RVT U1230 ( .A1(n470), .A2(n460), .Y(ab_13__15_) );
  AND2X1_RVT U1231 ( .A1(n470), .A2(n5), .Y(ab_13__14_) );
  AND2X1_RVT U1232 ( .A1(n470), .A2(n458), .Y(ab_13__13_) );
  AND2X1_RVT U1233 ( .A1(n470), .A2(n457), .Y(ab_13__12_) );
  AND2X1_RVT U1234 ( .A1(n470), .A2(n24), .Y(ab_13__11_) );
  AND2X1_RVT U1235 ( .A1(n470), .A2(n455), .Y(ab_13__10_) );
  AND2X1_RVT U1236 ( .A1(n470), .A2(n482), .Y(ab_13__0_) );
  AND2X1_RVT U1237 ( .A1(n469), .A2(n238), .Y(ab_12__9_) );
  AND2X1_RVT U1238 ( .A1(n469), .A2(n39), .Y(ab_12__8_) );
  AND2X1_RVT U1239 ( .A1(n469), .A2(n239), .Y(ab_12__7_) );
  AND2X1_RVT U1240 ( .A1(n469), .A2(n56), .Y(ab_12__6_) );
  AND2X1_RVT U1241 ( .A1(n469), .A2(n492), .Y(ab_12__5_) );
  AND2X1_RVT U1242 ( .A1(A[12]), .A2(n489), .Y(ab_12__4_) );
  AND2X1_RVT U1243 ( .A1(n469), .A2(n487), .Y(ab_12__3_) );
  AND2X1_RVT U1244 ( .A1(A[12]), .A2(n486), .Y(ab_12__2_) );
  AND2X1_RVT U1245 ( .A1(n469), .A2(n484), .Y(ab_12__1_) );
  AND2X1_RVT U1246 ( .A1(A[12]), .A2(n462), .Y(ab_12__19_) );
  AND2X1_RVT U1247 ( .A1(n469), .A2(n220), .Y(ab_12__18_) );
  AND2X1_RVT U1248 ( .A1(n469), .A2(n224), .Y(ab_12__17_) );
  AND2X1_RVT U1249 ( .A1(n469), .A2(n143), .Y(ab_12__16_) );
  AND2X1_RVT U1250 ( .A1(A[12]), .A2(n460), .Y(ab_12__15_) );
  AND2X1_RVT U1251 ( .A1(n469), .A2(n5), .Y(ab_12__14_) );
  AND2X1_RVT U1252 ( .A1(n469), .A2(n458), .Y(ab_12__13_) );
  AND2X1_RVT U1253 ( .A1(n469), .A2(n457), .Y(ab_12__12_) );
  AND2X1_RVT U1254 ( .A1(n469), .A2(n24), .Y(ab_12__11_) );
  AND2X1_RVT U1255 ( .A1(n469), .A2(n455), .Y(ab_12__10_) );
  AND2X1_RVT U1256 ( .A1(A[12]), .A2(n482), .Y(ab_12__0_) );
  AND2X1_RVT U1257 ( .A1(n467), .A2(n238), .Y(ab_11__9_) );
  AND2X1_RVT U1258 ( .A1(n468), .A2(n39), .Y(ab_11__8_) );
  AND2X1_RVT U1259 ( .A1(n467), .A2(n239), .Y(ab_11__7_) );
  AND2X1_RVT U1260 ( .A1(n468), .A2(n56), .Y(ab_11__6_) );
  AND2X1_RVT U1261 ( .A1(n467), .A2(n492), .Y(ab_11__5_) );
  AND2X1_RVT U1262 ( .A1(n468), .A2(n490), .Y(ab_11__4_) );
  AND2X1_RVT U1263 ( .A1(n467), .A2(n487), .Y(ab_11__3_) );
  AND2X1_RVT U1264 ( .A1(n468), .A2(n486), .Y(ab_11__2_) );
  AND2X1_RVT U1265 ( .A1(n467), .A2(n277), .Y(ab_11__20_) );
  AND2X1_RVT U1266 ( .A1(n468), .A2(n484), .Y(ab_11__1_) );
  AND2X1_RVT U1267 ( .A1(n467), .A2(n462), .Y(ab_11__19_) );
  AND2X1_RVT U1268 ( .A1(n468), .A2(n220), .Y(ab_11__18_) );
  AND2X1_RVT U1269 ( .A1(n467), .A2(n224), .Y(ab_11__17_) );
  AND2X1_RVT U1270 ( .A1(n468), .A2(n143), .Y(ab_11__16_) );
  AND2X1_RVT U1271 ( .A1(n467), .A2(n460), .Y(ab_11__15_) );
  AND2X1_RVT U1272 ( .A1(n468), .A2(n5), .Y(ab_11__14_) );
  AND2X1_RVT U1273 ( .A1(n467), .A2(n458), .Y(ab_11__13_) );
  AND2X1_RVT U1274 ( .A1(n468), .A2(n457), .Y(ab_11__12_) );
  AND2X1_RVT U1275 ( .A1(n467), .A2(n24), .Y(ab_11__11_) );
  AND2X1_RVT U1276 ( .A1(n468), .A2(n455), .Y(ab_11__10_) );
  AND2X1_RVT U1277 ( .A1(n467), .A2(n482), .Y(ab_11__0_) );
  AND2X1_RVT U1278 ( .A1(n465), .A2(n238), .Y(ab_10__9_) );
  AND2X1_RVT U1279 ( .A1(n466), .A2(n39), .Y(ab_10__8_) );
  AND2X1_RVT U1280 ( .A1(n465), .A2(n239), .Y(ab_10__7_) );
  AND2X1_RVT U1281 ( .A1(n466), .A2(n56), .Y(ab_10__6_) );
  AND2X1_RVT U1282 ( .A1(n465), .A2(n492), .Y(ab_10__5_) );
  AND2X1_RVT U1283 ( .A1(n466), .A2(n489), .Y(ab_10__4_) );
  AND2X1_RVT U1284 ( .A1(n465), .A2(n488), .Y(ab_10__3_) );
  AND2X1_RVT U1285 ( .A1(n466), .A2(n486), .Y(ab_10__2_) );
  AND2X1_RVT U1286 ( .A1(n465), .A2(n148), .Y(ab_10__21_) );
  AND2X1_RVT U1287 ( .A1(n466), .A2(n277), .Y(ab_10__20_) );
  AND2X1_RVT U1288 ( .A1(n465), .A2(n484), .Y(ab_10__1_) );
  AND2X1_RVT U1289 ( .A1(n466), .A2(n462), .Y(ab_10__19_) );
  AND2X1_RVT U1290 ( .A1(n465), .A2(n220), .Y(ab_10__18_) );
  AND2X1_RVT U1291 ( .A1(n466), .A2(n224), .Y(ab_10__17_) );
  AND2X1_RVT U1292 ( .A1(n465), .A2(n143), .Y(ab_10__16_) );
  AND2X1_RVT U1293 ( .A1(n466), .A2(n460), .Y(ab_10__15_) );
  AND2X1_RVT U1294 ( .A1(n465), .A2(n5), .Y(ab_10__14_) );
  AND2X1_RVT U1295 ( .A1(n466), .A2(n458), .Y(ab_10__13_) );
  AND2X1_RVT U1296 ( .A1(n465), .A2(n457), .Y(ab_10__12_) );
  AND2X1_RVT U1297 ( .A1(n466), .A2(n24), .Y(ab_10__11_) );
  AND2X1_RVT U1298 ( .A1(n465), .A2(n455), .Y(ab_10__10_) );
  AND2X1_RVT U1299 ( .A1(n466), .A2(n482), .Y(ab_10__0_) );
  AND2X1_RVT U1300 ( .A1(n57), .A2(B[8]), .Y(ab_0__8_) );
  AND2X1_RVT U1301 ( .A1(n381), .A2(n161), .Y(ab_0__7_) );
  AND2X1_RVT U1302 ( .A1(n381), .A2(n489), .Y(ab_0__4_) );
  AND2X1_RVT U1303 ( .A1(n325), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U1304 ( .A1(n325), .A2(n486), .Y(ab_0__2_) );
  AND2X1_RVT U1305 ( .A1(n57), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U1306 ( .A1(n57), .A2(B[16]), .Y(ab_0__16_) );
  AND2X1_RVT U1307 ( .A1(n57), .A2(B[14]), .Y(ab_0__14_) );
endmodule


module OSPE_0_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR3X2_RVT U1_31 ( .A1(A[31]), .A2(B[31]), .A3(carry[31]), .Y(SUM[31]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_0 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n44), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U8 ( .A1(n42), .A2(n47), .Y(N94) );
  AND2X1_RVT U13 ( .A1(n40), .A2(n46), .Y(N89) );
  AND2X1_RVT U19 ( .A1(n29), .A2(n44), .Y(N83) );
  AND2X1_RVT U25 ( .A1(n8), .A2(n44), .Y(N77) );
  AND2X1_RVT U26 ( .A1(n13), .A2(n44), .Y(N76) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n44), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n44), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n45), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n45), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n45), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n45), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n45), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n45), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n45), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n45), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n45), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n45), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n45), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n45), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n45), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n45), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n46), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n46), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n46), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n46), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n46), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n46), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n46), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n46), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n46), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n46), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n46), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n46), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n46), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n46), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n47), .Y(N44) );
  AND2X1_RVT U59 ( .A1(n12), .A2(n47), .Y(N43) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n49), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n49), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n49), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n48), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n49), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n49), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n49), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n49), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n49), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n49), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n49), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n49), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n48), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n48), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n48), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n48), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n48), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n48), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n48), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n48), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n48), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n48), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n48), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n48), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n48), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n48), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n49), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n49), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n49), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n49), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n49), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n47), .Y(N100) );
  OSPE_0_DW02_mult_0 mult_23 ( .A({ipA[31:5], n24, n33, ipA[2], n14, n39}), 
        .B({ipB[31:30], n41, n15, ipB[27], n31, n42, n34, n37, n36, n38, 
        ipB[20], n30, ipB[18], n2, n17, n21, n26, n9, n20, ipB[11], n1, 
        ipB[9:0]}), .PRODUCT_31_(N35), .PRODUCT_30_(N34), .PRODUCT_29_(N33), 
        .PRODUCT_28_(N32), .PRODUCT_27_(N31), .PRODUCT_26_(N30), .PRODUCT_25_(
        N29), .PRODUCT_24_(N28), .PRODUCT_23_(N27), .PRODUCT_22_(N26), 
        .PRODUCT_21_(N25), .PRODUCT_20_(N24), .PRODUCT_19_(N23), .PRODUCT_18_(
        N22), .PRODUCT_17_(N21), .PRODUCT_16_(N20), .PRODUCT_15_(N19), 
        .PRODUCT_14_(N18), .PRODUCT_13_(N17), .PRODUCT_12_(N16), .PRODUCT_11_(
        N15), .PRODUCT_10_(N14), .PRODUCT_9_(N13), .PRODUCT_8_(N12), 
        .PRODUCT_7_(N11), .PRODUCT_6_(N10), .PRODUCT_5_(N9), .PRODUCT_4_(N8), 
        .PRODUCT_3_(N7), .PRODUCT_2_(N6), .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_0_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX2_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  NBUFFX2_RVT U4 ( .A(ipB[10]), .Y(n1) );
  NBUFFX2_RVT U5 ( .A(ipB[17]), .Y(n2) );
  DELLN3X2_RVT U6 ( .A(n17), .Y(n3) );
  AND2X4_RVT U7 ( .A1(ipA[5]), .A2(n47), .Y(N42) );
  DELLN3X2_RVT U9 ( .A(n38), .Y(n4) );
  DELLN3X2_RVT U10 ( .A(n14), .Y(n5) );
  AND2X4_RVT U11 ( .A1(n5), .A2(n47), .Y(N38) );
  IBUFFX2_RVT U12 ( .A(n3), .Y(n6) );
  INVX1_RVT U14 ( .A(n6), .Y(n7) );
  DELLN3X2_RVT U15 ( .A(ipB[8]), .Y(n8) );
  NBUFFX2_RVT U16 ( .A(ipB[13]), .Y(n9) );
  AND2X1_RVT U17 ( .A1(n22), .A2(n46), .Y(N91) );
  AND2X1_RVT U18 ( .A1(n27), .A2(n47), .Y(N92) );
  AND2X1_RVT U20 ( .A1(n32), .A2(n47), .Y(N37) );
  AND2X1_RVT U21 ( .A1(ipA[2]), .A2(n47), .Y(N39) );
  AND2X1_RVT U22 ( .A1(n18), .A2(n44), .Y(N86) );
  AND2X1_RVT U23 ( .A1(n35), .A2(n47), .Y(N87) );
  AND2X1_RVT U24 ( .A1(n10), .A2(n47), .Y(N88) );
  AND2X1_RVT U27 ( .A1(n28), .A2(n47), .Y(N41) );
  AND2X1_RVT U60 ( .A1(n19), .A2(n44), .Y(N75) );
  AND2X1_RVT U61 ( .A1(n11), .A2(n44), .Y(N78) );
  AND2X1_RVT U62 ( .A1(n16), .A2(n44), .Y(N80) );
  AND2X1_RVT U63 ( .A1(n25), .A2(n44), .Y(N81) );
  AND2X1_RVT U64 ( .A1(n23), .A2(n44), .Y(N84) );
  AND2X4_RVT U65 ( .A1(n7), .A2(n44), .Y(N85) );
  DELLN3X2_RVT U66 ( .A(n30), .Y(n10) );
  DELLN3X2_RVT U99 ( .A(ipB[9]), .Y(n11) );
  AND2X4_RVT U100 ( .A1(n1), .A2(n44), .Y(N79) );
  DELLN3X2_RVT U101 ( .A(ipA[6]), .Y(n12) );
  DELLN3X2_RVT U102 ( .A(ipB[7]), .Y(n13) );
  NBUFFX2_RVT U103 ( .A(ipA[1]), .Y(n14) );
  AND2X1_RVT U104 ( .A1(rstnPsum), .A2(opC_wire[31]), .Y(N133) );
  NBUFFX2_RVT U105 ( .A(ipB[28]), .Y(n15) );
  DELLN3X2_RVT U106 ( .A(ipB[11]), .Y(n16) );
  NBUFFX2_RVT U107 ( .A(ipB[16]), .Y(n17) );
  DELLN3X2_RVT U108 ( .A(n2), .Y(n18) );
  DELLN3X2_RVT U109 ( .A(ipB[6]), .Y(n19) );
  AND2X4_RVT U110 ( .A1(n4), .A2(n47), .Y(N90) );
  AND2X4_RVT U111 ( .A1(n9), .A2(n44), .Y(N82) );
  NBUFFX2_RVT U112 ( .A(ipB[12]), .Y(n20) );
  NBUFFX2_RVT U113 ( .A(ipB[15]), .Y(n21) );
  DELLN3X2_RVT U114 ( .A(n36), .Y(n22) );
  AND2X4_RVT U115 ( .A1(ipB[27]), .A2(n47), .Y(N96) );
  DELLN3X2_RVT U116 ( .A(n21), .Y(n23) );
  AND2X4_RVT U117 ( .A1(n33), .A2(n47), .Y(N40) );
  NBUFFX2_RVT U118 ( .A(ipA[4]), .Y(n24) );
  DELLN3X2_RVT U119 ( .A(n20), .Y(n25) );
  NBUFFX2_RVT U120 ( .A(ipB[14]), .Y(n26) );
  NBUFFX2_RVT U121 ( .A(ipB[19]), .Y(n30) );
  DELLN3X2_RVT U122 ( .A(n37), .Y(n27) );
  DELLN3X2_RVT U123 ( .A(n24), .Y(n28) );
  DELLN3X2_RVT U124 ( .A(n26), .Y(n29) );
  NBUFFX2_RVT U125 ( .A(ipB[26]), .Y(n31) );
  DELLN3X2_RVT U126 ( .A(n39), .Y(n32) );
  NBUFFX2_RVT U127 ( .A(ipA[3]), .Y(n33) );
  NBUFFX2_RVT U128 ( .A(ipB[24]), .Y(n34) );
  DELLN3X2_RVT U129 ( .A(ipB[18]), .Y(n35) );
  AND2X4_RVT U130 ( .A1(n34), .A2(n45), .Y(N93) );
  NBUFFX2_RVT U131 ( .A(ipB[22]), .Y(n36) );
  NBUFFX2_RVT U132 ( .A(ipB[23]), .Y(n37) );
  NBUFFX2_RVT U133 ( .A(ipB[21]), .Y(n38) );
  NBUFFX2_RVT U134 ( .A(ipA[0]), .Y(n39) );
  DELLN3X2_RVT U135 ( .A(ipB[20]), .Y(n40) );
  DELLN3X2_RVT U136 ( .A(n41), .Y(n43) );
  AND2X4_RVT U137 ( .A1(n15), .A2(n47), .Y(N97) );
  AND2X4_RVT U138 ( .A1(n31), .A2(n44), .Y(N95) );
  NBUFFX2_RVT U139 ( .A(rstnPipe), .Y(n44) );
  NBUFFX2_RVT U140 ( .A(rstnPipe), .Y(n46) );
  NBUFFX2_RVT U141 ( .A(rstnPipe), .Y(n45) );
  NBUFFX2_RVT U142 ( .A(rstnPipe), .Y(n47) );
  AND2X1_RVT U143 ( .A1(n43), .A2(n45), .Y(N98) );
  NBUFFX2_RVT U144 ( .A(rstnPsum), .Y(n48) );
  NBUFFX2_RVT U145 ( .A(rstnPsum), .Y(n49) );
  NBUFFX2_RVT U146 ( .A(ipB[29]), .Y(n41) );
  NBUFFX2_RVT U147 ( .A(ipB[25]), .Y(n42) );
endmodule


module OSPE_15_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR2X1_RVT U16 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U17 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U18 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U19 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U20 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U21 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U22 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  NBUFFX2_RVT U23 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U25 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_15_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_15 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n1), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n4), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n1), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n4), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n1), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n4), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n4), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n4), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n4), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n4), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_15_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_15_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_14_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U5 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U6 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U7 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U8 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U9 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U10 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U11 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U12 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U13 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U14 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U15 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U16 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U17 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U18 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U19 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U20 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U21 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  XOR2X1_RVT U22 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U23 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U24 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR2X1_RVT U25 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U27 ( .A(A[1]), .Y(n38) );
  NBUFFX2_RVT U28 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U29 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U30 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U31 ( .A(A[3]), .Y(n42) );
  XOR2X1_RVT U32 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U33 ( .A(A[0]), .Y(n36) );
  NBUFFX2_RVT U34 ( .A(A[1]), .Y(n39) );
  XOR2X1_RVT U35 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U36 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U37 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U38 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U39 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n41) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n63) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n75) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n73) );
  NBUFFX2_RVT U44 ( .A(B[7]), .Y(n71) );
  NBUFFX2_RVT U45 ( .A(A[9]), .Y(n55) );
  NBUFFX2_RVT U46 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U47 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U48 ( .A(B[6]), .Y(n69) );
  NBUFFX2_RVT U49 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U50 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U51 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U52 ( .A(B[5]), .Y(n66) );
  NBUFFX2_RVT U53 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U54 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U55 ( .A(B[4]), .Y(n65) );
  NBUFFX2_RVT U56 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U57 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U58 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U59 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U60 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U61 ( .A(A[6]), .Y(n48) );
  NBUFFX2_RVT U62 ( .A(A[7]), .Y(n51) );
  NBUFFX2_RVT U63 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U64 ( .A(B[5]), .Y(n67) );
  NBUFFX2_RVT U65 ( .A(A[8]), .Y(n53) );
  NBUFFX2_RVT U66 ( .A(A[8]), .Y(n52) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n43) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n57) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n45) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n59) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n47) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n61) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n49) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  NBUFFX2_RVT U116 ( .A(B[19]), .Y(n14) );
  NBUFFX2_RVT U117 ( .A(B[20]), .Y(n15) );
  NBUFFX2_RVT U118 ( .A(B[21]), .Y(n16) );
  NBUFFX2_RVT U119 ( .A(B[22]), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(B[23]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[10]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[11]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[12]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[13]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[14]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[15]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[16]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[17]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[18]), .Y(n28) );
  NBUFFX2_RVT U131 ( .A(A[19]), .Y(n29) );
  INVX0_RVT U132 ( .A(A[20]), .Y(n30) );
  INVX0_RVT U133 ( .A(n30), .Y(n31) );
  INVX0_RVT U134 ( .A(A[21]), .Y(n32) );
  INVX0_RVT U135 ( .A(n32), .Y(n33) );
  AND2X1_RVT U136 ( .A1(n74), .A2(n55), .Y(ab_9__9_) );
  AND2X1_RVT U137 ( .A1(n72), .A2(n55), .Y(ab_9__8_) );
  AND2X1_RVT U138 ( .A1(n70), .A2(n55), .Y(ab_9__7_) );
  AND2X1_RVT U139 ( .A1(n68), .A2(n55), .Y(ab_9__6_) );
  AND2X1_RVT U140 ( .A1(n66), .A2(n55), .Y(ab_9__5_) );
  AND2X1_RVT U141 ( .A1(n64), .A2(n55), .Y(ab_9__4_) );
  AND2X1_RVT U142 ( .A1(n63), .A2(n55), .Y(ab_9__3_) );
  AND2X1_RVT U143 ( .A1(n61), .A2(n55), .Y(ab_9__2_) );
  AND2X1_RVT U144 ( .A1(n17), .A2(n55), .Y(ab_9__22_) );
  AND2X1_RVT U145 ( .A1(n16), .A2(n55), .Y(ab_9__21_) );
  AND2X1_RVT U146 ( .A1(n15), .A2(n55), .Y(ab_9__20_) );
  AND2X1_RVT U147 ( .A1(n59), .A2(n54), .Y(ab_9__1_) );
  AND2X1_RVT U148 ( .A1(n14), .A2(n54), .Y(ab_9__19_) );
  AND2X1_RVT U149 ( .A1(n13), .A2(n54), .Y(ab_9__18_) );
  AND2X1_RVT U150 ( .A1(B[17]), .A2(n54), .Y(ab_9__17_) );
  AND2X1_RVT U151 ( .A1(n11), .A2(n54), .Y(ab_9__16_) );
  AND2X1_RVT U152 ( .A1(n10), .A2(n54), .Y(ab_9__15_) );
  AND2X1_RVT U153 ( .A1(n9), .A2(n54), .Y(ab_9__14_) );
  AND2X1_RVT U154 ( .A1(B[13]), .A2(n54), .Y(ab_9__13_) );
  AND2X1_RVT U155 ( .A1(n7), .A2(n54), .Y(ab_9__12_) );
  AND2X1_RVT U156 ( .A1(n5), .A2(n54), .Y(ab_9__11_) );
  AND2X1_RVT U157 ( .A1(n3), .A2(n54), .Y(ab_9__10_) );
  AND2X1_RVT U158 ( .A1(n56), .A2(n54), .Y(ab_9__0_) );
  AND2X1_RVT U159 ( .A1(n53), .A2(n74), .Y(ab_8__9_) );
  AND2X1_RVT U160 ( .A1(n53), .A2(n72), .Y(ab_8__8_) );
  AND2X1_RVT U161 ( .A1(n53), .A2(n70), .Y(ab_8__7_) );
  AND2X1_RVT U162 ( .A1(n53), .A2(n68), .Y(ab_8__6_) );
  AND2X1_RVT U163 ( .A1(n53), .A2(n66), .Y(ab_8__5_) );
  AND2X1_RVT U164 ( .A1(n53), .A2(n64), .Y(ab_8__4_) );
  AND2X1_RVT U165 ( .A1(n53), .A2(n63), .Y(ab_8__3_) );
  AND2X1_RVT U166 ( .A1(n53), .A2(n61), .Y(ab_8__2_) );
  AND2X1_RVT U167 ( .A1(n53), .A2(n18), .Y(ab_8__23_) );
  AND2X1_RVT U168 ( .A1(n53), .A2(n17), .Y(ab_8__22_) );
  AND2X1_RVT U169 ( .A1(n53), .A2(n16), .Y(ab_8__21_) );
  AND2X1_RVT U170 ( .A1(n53), .A2(n15), .Y(ab_8__20_) );
  AND2X1_RVT U171 ( .A1(n52), .A2(n59), .Y(ab_8__1_) );
  AND2X1_RVT U172 ( .A1(n52), .A2(n14), .Y(ab_8__19_) );
  AND2X1_RVT U173 ( .A1(n52), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U174 ( .A1(n52), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U175 ( .A1(n52), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U176 ( .A1(n52), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U177 ( .A1(n52), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U178 ( .A1(n52), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U179 ( .A1(n52), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U180 ( .A1(n52), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U181 ( .A1(n52), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U182 ( .A1(n52), .A2(n56), .Y(ab_8__0_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n74), .Y(ab_7__9_) );
  AND2X1_RVT U184 ( .A1(n51), .A2(n72), .Y(ab_7__8_) );
  AND2X1_RVT U185 ( .A1(n51), .A2(n70), .Y(ab_7__7_) );
  AND2X1_RVT U186 ( .A1(n51), .A2(n68), .Y(ab_7__6_) );
  AND2X1_RVT U187 ( .A1(n51), .A2(n66), .Y(ab_7__5_) );
  AND2X1_RVT U188 ( .A1(n51), .A2(n64), .Y(ab_7__4_) );
  AND2X1_RVT U189 ( .A1(n51), .A2(n63), .Y(ab_7__3_) );
  AND2X1_RVT U190 ( .A1(n51), .A2(n61), .Y(ab_7__2_) );
  AND2X1_RVT U191 ( .A1(n51), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U192 ( .A1(n51), .A2(n18), .Y(ab_7__23_) );
  AND2X1_RVT U193 ( .A1(n51), .A2(n17), .Y(ab_7__22_) );
  AND2X1_RVT U194 ( .A1(n51), .A2(n16), .Y(ab_7__21_) );
  AND2X1_RVT U195 ( .A1(n51), .A2(n15), .Y(ab_7__20_) );
  AND2X1_RVT U196 ( .A1(n50), .A2(n59), .Y(ab_7__1_) );
  AND2X1_RVT U197 ( .A1(n50), .A2(n14), .Y(ab_7__19_) );
  AND2X1_RVT U198 ( .A1(n50), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U199 ( .A1(n50), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U200 ( .A1(n50), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U201 ( .A1(n50), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U202 ( .A1(n50), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U203 ( .A1(n50), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U204 ( .A1(n50), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U205 ( .A1(n50), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U206 ( .A1(n50), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U207 ( .A1(n50), .A2(n56), .Y(ab_7__0_) );
  AND2X1_RVT U208 ( .A1(n49), .A2(n74), .Y(ab_6__9_) );
  AND2X1_RVT U209 ( .A1(n49), .A2(n72), .Y(ab_6__8_) );
  AND2X1_RVT U210 ( .A1(n48), .A2(n70), .Y(ab_6__7_) );
  AND2X1_RVT U211 ( .A1(n48), .A2(n68), .Y(ab_6__6_) );
  AND2X1_RVT U212 ( .A1(n48), .A2(n66), .Y(ab_6__5_) );
  AND2X1_RVT U213 ( .A1(n48), .A2(n64), .Y(ab_6__4_) );
  AND2X1_RVT U214 ( .A1(n48), .A2(n63), .Y(ab_6__3_) );
  AND2X1_RVT U215 ( .A1(n48), .A2(n61), .Y(ab_6__2_) );
  AND2X1_RVT U216 ( .A1(n48), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U217 ( .A1(n48), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U218 ( .A1(n48), .A2(n18), .Y(ab_6__23_) );
  AND2X1_RVT U219 ( .A1(n48), .A2(n17), .Y(ab_6__22_) );
  AND2X1_RVT U220 ( .A1(n48), .A2(n16), .Y(ab_6__21_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n15), .Y(ab_6__20_) );
  AND2X1_RVT U222 ( .A1(n49), .A2(n59), .Y(ab_6__1_) );
  AND2X1_RVT U223 ( .A1(n49), .A2(n14), .Y(ab_6__19_) );
  AND2X1_RVT U224 ( .A1(n49), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U225 ( .A1(n49), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U226 ( .A1(n49), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U227 ( .A1(n49), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U228 ( .A1(n49), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U229 ( .A1(n49), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U230 ( .A1(n49), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U231 ( .A1(n49), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U232 ( .A1(n49), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U233 ( .A1(n49), .A2(n56), .Y(ab_6__0_) );
  AND2X1_RVT U234 ( .A1(n47), .A2(n74), .Y(ab_5__9_) );
  AND2X1_RVT U235 ( .A1(n47), .A2(n72), .Y(ab_5__8_) );
  AND2X1_RVT U236 ( .A1(n47), .A2(n70), .Y(ab_5__7_) );
  AND2X1_RVT U237 ( .A1(n46), .A2(n68), .Y(ab_5__6_) );
  AND2X1_RVT U238 ( .A1(n46), .A2(n66), .Y(ab_5__5_) );
  AND2X1_RVT U239 ( .A1(n46), .A2(n64), .Y(ab_5__4_) );
  AND2X1_RVT U240 ( .A1(n46), .A2(n63), .Y(ab_5__3_) );
  AND2X1_RVT U241 ( .A1(n46), .A2(n61), .Y(ab_5__2_) );
  AND2X1_RVT U242 ( .A1(n46), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U243 ( .A1(n46), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U244 ( .A1(n46), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U245 ( .A1(n46), .A2(n18), .Y(ab_5__23_) );
  AND2X1_RVT U246 ( .A1(n46), .A2(n17), .Y(ab_5__22_) );
  AND2X1_RVT U247 ( .A1(n46), .A2(n16), .Y(ab_5__21_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n15), .Y(ab_5__20_) );
  AND2X1_RVT U249 ( .A1(n47), .A2(n59), .Y(ab_5__1_) );
  AND2X1_RVT U250 ( .A1(n47), .A2(n14), .Y(ab_5__19_) );
  AND2X1_RVT U251 ( .A1(n47), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U252 ( .A1(n47), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U253 ( .A1(n47), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U254 ( .A1(n47), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U255 ( .A1(n47), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U256 ( .A1(n47), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U257 ( .A1(n47), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U258 ( .A1(n47), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U259 ( .A1(n47), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U260 ( .A1(n47), .A2(n56), .Y(ab_5__0_) );
  AND2X1_RVT U261 ( .A1(n45), .A2(n74), .Y(ab_4__9_) );
  AND2X1_RVT U262 ( .A1(n45), .A2(n72), .Y(ab_4__8_) );
  AND2X1_RVT U263 ( .A1(n45), .A2(n70), .Y(ab_4__7_) );
  AND2X1_RVT U264 ( .A1(n45), .A2(n68), .Y(ab_4__6_) );
  AND2X1_RVT U265 ( .A1(n44), .A2(n66), .Y(ab_4__5_) );
  AND2X1_RVT U266 ( .A1(n44), .A2(n64), .Y(ab_4__4_) );
  AND2X1_RVT U267 ( .A1(n44), .A2(n63), .Y(ab_4__3_) );
  AND2X1_RVT U268 ( .A1(n44), .A2(n61), .Y(ab_4__2_) );
  AND2X1_RVT U269 ( .A1(n44), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U270 ( .A1(n44), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U271 ( .A1(n44), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U272 ( .A1(n44), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U273 ( .A1(n44), .A2(n18), .Y(ab_4__23_) );
  AND2X1_RVT U274 ( .A1(n44), .A2(n17), .Y(ab_4__22_) );
  AND2X1_RVT U275 ( .A1(n44), .A2(n16), .Y(ab_4__21_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n15), .Y(ab_4__20_) );
  AND2X1_RVT U277 ( .A1(n45), .A2(n59), .Y(ab_4__1_) );
  AND2X1_RVT U278 ( .A1(n45), .A2(n14), .Y(ab_4__19_) );
  AND2X1_RVT U279 ( .A1(n45), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U280 ( .A1(n45), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U281 ( .A1(n45), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U282 ( .A1(n45), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U283 ( .A1(n45), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U284 ( .A1(n45), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U285 ( .A1(n45), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U286 ( .A1(n45), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U287 ( .A1(n45), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U288 ( .A1(n45), .A2(n56), .Y(ab_4__0_) );
  AND2X1_RVT U289 ( .A1(n43), .A2(n74), .Y(ab_3__9_) );
  AND2X1_RVT U290 ( .A1(n43), .A2(n72), .Y(ab_3__8_) );
  AND2X1_RVT U291 ( .A1(n43), .A2(n70), .Y(ab_3__7_) );
  AND2X1_RVT U292 ( .A1(n43), .A2(n68), .Y(ab_3__6_) );
  AND2X1_RVT U293 ( .A1(n43), .A2(n66), .Y(ab_3__5_) );
  AND2X1_RVT U294 ( .A1(n42), .A2(n64), .Y(ab_3__4_) );
  AND2X1_RVT U295 ( .A1(n42), .A2(n63), .Y(ab_3__3_) );
  AND2X1_RVT U296 ( .A1(n42), .A2(n61), .Y(ab_3__2_) );
  AND2X1_RVT U297 ( .A1(n42), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U298 ( .A1(n42), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U299 ( .A1(n42), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U300 ( .A1(n42), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U301 ( .A1(n42), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U302 ( .A1(n42), .A2(n18), .Y(ab_3__23_) );
  AND2X1_RVT U303 ( .A1(n42), .A2(n17), .Y(ab_3__22_) );
  AND2X1_RVT U304 ( .A1(n42), .A2(n16), .Y(ab_3__21_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n15), .Y(ab_3__20_) );
  AND2X1_RVT U306 ( .A1(n43), .A2(n59), .Y(ab_3__1_) );
  AND2X1_RVT U307 ( .A1(n43), .A2(n14), .Y(ab_3__19_) );
  AND2X1_RVT U308 ( .A1(n43), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U309 ( .A1(n43), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U310 ( .A1(n43), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U311 ( .A1(n43), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U312 ( .A1(n43), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U313 ( .A1(n43), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U314 ( .A1(n43), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U315 ( .A1(n43), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U316 ( .A1(n43), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U317 ( .A1(n43), .A2(n56), .Y(ab_3__0_) );
  AND2X1_RVT U318 ( .A1(A[31]), .A2(n56), .Y(ab_31__0_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n59), .Y(ab_30__1_) );
  AND2X1_RVT U320 ( .A1(A[30]), .A2(n56), .Y(ab_30__0_) );
  AND2X1_RVT U321 ( .A1(n41), .A2(n74), .Y(ab_2__9_) );
  AND2X1_RVT U322 ( .A1(n41), .A2(n72), .Y(ab_2__8_) );
  AND2X1_RVT U323 ( .A1(n41), .A2(n70), .Y(ab_2__7_) );
  AND2X1_RVT U324 ( .A1(n41), .A2(n68), .Y(ab_2__6_) );
  AND2X1_RVT U325 ( .A1(n41), .A2(n66), .Y(ab_2__5_) );
  AND2X1_RVT U326 ( .A1(n41), .A2(n64), .Y(ab_2__4_) );
  AND2X1_RVT U327 ( .A1(n41), .A2(n63), .Y(ab_2__3_) );
  AND2X1_RVT U328 ( .A1(n40), .A2(n61), .Y(ab_2__2_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U330 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U331 ( .A1(n41), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U332 ( .A1(n40), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U333 ( .A1(n40), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U334 ( .A1(n40), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U335 ( .A1(A[2]), .A2(n18), .Y(ab_2__23_) );
  AND2X1_RVT U336 ( .A1(n41), .A2(n17), .Y(ab_2__22_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n16), .Y(ab_2__21_) );
  AND2X1_RVT U338 ( .A1(A[2]), .A2(n15), .Y(ab_2__20_) );
  AND2X1_RVT U339 ( .A1(n40), .A2(n59), .Y(ab_2__1_) );
  AND2X1_RVT U340 ( .A1(n40), .A2(n14), .Y(ab_2__19_) );
  AND2X1_RVT U341 ( .A1(n40), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U342 ( .A1(n40), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U343 ( .A1(n40), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U344 ( .A1(n40), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U345 ( .A1(n40), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U346 ( .A1(n40), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U347 ( .A1(n40), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U348 ( .A1(n40), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U349 ( .A1(n40), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U350 ( .A1(n40), .A2(n56), .Y(ab_2__0_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n61), .Y(ab_29__2_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n59), .Y(ab_29__1_) );
  AND2X1_RVT U353 ( .A1(A[29]), .A2(n56), .Y(ab_29__0_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n63), .Y(ab_28__3_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n61), .Y(ab_28__2_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n59), .Y(ab_28__1_) );
  AND2X1_RVT U357 ( .A1(A[28]), .A2(n56), .Y(ab_28__0_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n64), .Y(ab_27__4_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n63), .Y(ab_27__3_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n61), .Y(ab_27__2_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n59), .Y(ab_27__1_) );
  AND2X1_RVT U362 ( .A1(A[27]), .A2(n56), .Y(ab_27__0_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n66), .Y(ab_26__5_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n64), .Y(ab_26__4_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n63), .Y(ab_26__3_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n61), .Y(ab_26__2_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n59), .Y(ab_26__1_) );
  AND2X1_RVT U368 ( .A1(A[26]), .A2(n57), .Y(ab_26__0_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n68), .Y(ab_25__6_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n66), .Y(ab_25__5_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n64), .Y(ab_25__4_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n63), .Y(ab_25__3_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n61), .Y(ab_25__2_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n58), .Y(ab_25__1_) );
  AND2X1_RVT U375 ( .A1(A[25]), .A2(n57), .Y(ab_25__0_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n70), .Y(ab_24__7_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n68), .Y(ab_24__6_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n66), .Y(ab_24__5_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n64), .Y(ab_24__4_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n63), .Y(ab_24__3_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n60), .Y(ab_24__2_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n58), .Y(ab_24__1_) );
  AND2X1_RVT U383 ( .A1(A[24]), .A2(n57), .Y(ab_24__0_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n72), .Y(ab_23__8_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n70), .Y(ab_23__7_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n68), .Y(ab_23__6_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n66), .Y(ab_23__5_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n64), .Y(ab_23__4_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n62), .Y(ab_23__3_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n60), .Y(ab_23__2_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n58), .Y(ab_23__1_) );
  AND2X1_RVT U392 ( .A1(A[23]), .A2(n57), .Y(ab_23__0_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n74), .Y(ab_22__9_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n72), .Y(ab_22__8_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n70), .Y(ab_22__7_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n68), .Y(ab_22__6_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n66), .Y(ab_22__5_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n65), .Y(ab_22__4_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n62), .Y(ab_22__3_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n60), .Y(ab_22__2_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n58), .Y(ab_22__1_) );
  AND2X1_RVT U402 ( .A1(A[22]), .A2(n57), .Y(ab_22__0_) );
  AND2X1_RVT U403 ( .A1(A[21]), .A2(n74), .Y(ab_21__9_) );
  AND2X1_RVT U404 ( .A1(n33), .A2(n72), .Y(ab_21__8_) );
  AND2X1_RVT U405 ( .A1(n33), .A2(n70), .Y(ab_21__7_) );
  AND2X1_RVT U406 ( .A1(n33), .A2(n68), .Y(ab_21__6_) );
  AND2X1_RVT U407 ( .A1(n33), .A2(n67), .Y(ab_21__5_) );
  AND2X1_RVT U408 ( .A1(n33), .A2(n65), .Y(ab_21__4_) );
  AND2X1_RVT U409 ( .A1(n33), .A2(n62), .Y(ab_21__3_) );
  AND2X1_RVT U410 ( .A1(n33), .A2(n60), .Y(ab_21__2_) );
  AND2X1_RVT U411 ( .A1(n33), .A2(n58), .Y(ab_21__1_) );
  AND2X1_RVT U412 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U413 ( .A1(n33), .A2(n57), .Y(ab_21__0_) );
  AND2X1_RVT U414 ( .A1(n31), .A2(n74), .Y(ab_20__9_) );
  AND2X1_RVT U415 ( .A1(n31), .A2(n72), .Y(ab_20__8_) );
  AND2X1_RVT U416 ( .A1(n31), .A2(n70), .Y(ab_20__7_) );
  AND2X1_RVT U417 ( .A1(n31), .A2(n69), .Y(ab_20__6_) );
  AND2X1_RVT U418 ( .A1(n31), .A2(n67), .Y(ab_20__5_) );
  AND2X1_RVT U419 ( .A1(n31), .A2(n65), .Y(ab_20__4_) );
  AND2X1_RVT U420 ( .A1(n31), .A2(n62), .Y(ab_20__3_) );
  AND2X1_RVT U421 ( .A1(n31), .A2(n60), .Y(ab_20__2_) );
  AND2X1_RVT U422 ( .A1(n31), .A2(n58), .Y(ab_20__1_) );
  AND2X1_RVT U423 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U424 ( .A1(n31), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U425 ( .A1(n31), .A2(n57), .Y(ab_20__0_) );
  AND2X1_RVT U426 ( .A1(n39), .A2(n74), .Y(ab_1__9_) );
  AND2X1_RVT U427 ( .A1(n39), .A2(n72), .Y(ab_1__8_) );
  AND2X1_RVT U428 ( .A1(n39), .A2(n71), .Y(ab_1__7_) );
  AND2X1_RVT U429 ( .A1(n39), .A2(n69), .Y(ab_1__6_) );
  AND2X1_RVT U430 ( .A1(n39), .A2(n67), .Y(ab_1__5_) );
  AND2X1_RVT U431 ( .A1(n39), .A2(n65), .Y(ab_1__4_) );
  AND2X1_RVT U432 ( .A1(n39), .A2(n62), .Y(ab_1__3_) );
  AND2X1_RVT U433 ( .A1(n38), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U434 ( .A1(n38), .A2(n60), .Y(ab_1__2_) );
  AND2X1_RVT U435 ( .A1(n38), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U436 ( .A1(n38), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U437 ( .A1(n38), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U438 ( .A1(n38), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U439 ( .A1(n38), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U440 ( .A1(n38), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U441 ( .A1(n38), .A2(n18), .Y(ab_1__23_) );
  AND2X1_RVT U442 ( .A1(n38), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U443 ( .A1(n38), .A2(n16), .Y(ab_1__21_) );
  AND2X1_RVT U444 ( .A1(n38), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U445 ( .A1(n37), .A2(n58), .Y(ab_1__1_) );
  AND2X1_RVT U446 ( .A1(n37), .A2(n14), .Y(ab_1__19_) );
  AND2X1_RVT U447 ( .A1(n37), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U448 ( .A1(n37), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U449 ( .A1(n37), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U450 ( .A1(n37), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U451 ( .A1(n37), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U452 ( .A1(n37), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U453 ( .A1(n37), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U454 ( .A1(n37), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U455 ( .A1(n37), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U456 ( .A1(n37), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U457 ( .A1(n29), .A2(n74), .Y(ab_19__9_) );
  AND2X1_RVT U458 ( .A1(n29), .A2(n73), .Y(ab_19__8_) );
  AND2X1_RVT U459 ( .A1(n29), .A2(n71), .Y(ab_19__7_) );
  AND2X1_RVT U460 ( .A1(n29), .A2(n69), .Y(ab_19__6_) );
  AND2X1_RVT U461 ( .A1(n29), .A2(n67), .Y(ab_19__5_) );
  AND2X1_RVT U462 ( .A1(n29), .A2(n65), .Y(ab_19__4_) );
  AND2X1_RVT U463 ( .A1(n29), .A2(n62), .Y(ab_19__3_) );
  AND2X1_RVT U464 ( .A1(n29), .A2(n60), .Y(ab_19__2_) );
  AND2X1_RVT U465 ( .A1(n29), .A2(n58), .Y(ab_19__1_) );
  AND2X1_RVT U466 ( .A1(n29), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U467 ( .A1(n29), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U468 ( .A1(n29), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U469 ( .A1(A[19]), .A2(n57), .Y(ab_19__0_) );
  AND2X1_RVT U470 ( .A1(n28), .A2(n75), .Y(ab_18__9_) );
  AND2X1_RVT U471 ( .A1(n28), .A2(n73), .Y(ab_18__8_) );
  AND2X1_RVT U472 ( .A1(n28), .A2(n71), .Y(ab_18__7_) );
  AND2X1_RVT U473 ( .A1(n28), .A2(n69), .Y(ab_18__6_) );
  AND2X1_RVT U474 ( .A1(n28), .A2(n67), .Y(ab_18__5_) );
  AND2X1_RVT U475 ( .A1(n28), .A2(n65), .Y(ab_18__4_) );
  AND2X1_RVT U476 ( .A1(n28), .A2(n62), .Y(ab_18__3_) );
  AND2X1_RVT U477 ( .A1(n28), .A2(n60), .Y(ab_18__2_) );
  AND2X1_RVT U478 ( .A1(A[18]), .A2(n58), .Y(ab_18__1_) );
  AND2X1_RVT U479 ( .A1(n28), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U480 ( .A1(n28), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U481 ( .A1(n28), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U482 ( .A1(n28), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U483 ( .A1(n28), .A2(n57), .Y(ab_18__0_) );
  AND2X1_RVT U484 ( .A1(n27), .A2(n75), .Y(ab_17__9_) );
  AND2X1_RVT U485 ( .A1(n27), .A2(n73), .Y(ab_17__8_) );
  AND2X1_RVT U486 ( .A1(n27), .A2(n71), .Y(ab_17__7_) );
  AND2X1_RVT U487 ( .A1(n27), .A2(n69), .Y(ab_17__6_) );
  AND2X1_RVT U488 ( .A1(n27), .A2(n67), .Y(ab_17__5_) );
  AND2X1_RVT U489 ( .A1(n27), .A2(n65), .Y(ab_17__4_) );
  AND2X1_RVT U490 ( .A1(n27), .A2(n62), .Y(ab_17__3_) );
  AND2X1_RVT U491 ( .A1(n27), .A2(n60), .Y(ab_17__2_) );
  AND2X1_RVT U492 ( .A1(A[17]), .A2(n58), .Y(ab_17__1_) );
  AND2X1_RVT U493 ( .A1(n27), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U494 ( .A1(n27), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U495 ( .A1(n27), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U496 ( .A1(n27), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U497 ( .A1(n27), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U498 ( .A1(A[17]), .A2(n57), .Y(ab_17__0_) );
  AND2X1_RVT U499 ( .A1(n26), .A2(n75), .Y(ab_16__9_) );
  AND2X1_RVT U500 ( .A1(n26), .A2(n73), .Y(ab_16__8_) );
  AND2X1_RVT U501 ( .A1(n26), .A2(n71), .Y(ab_16__7_) );
  AND2X1_RVT U502 ( .A1(n26), .A2(n69), .Y(ab_16__6_) );
  AND2X1_RVT U503 ( .A1(n26), .A2(n67), .Y(ab_16__5_) );
  AND2X1_RVT U504 ( .A1(n26), .A2(n65), .Y(ab_16__4_) );
  AND2X1_RVT U505 ( .A1(A[16]), .A2(n62), .Y(ab_16__3_) );
  AND2X1_RVT U506 ( .A1(n26), .A2(n60), .Y(ab_16__2_) );
  AND2X1_RVT U507 ( .A1(A[16]), .A2(n58), .Y(ab_16__1_) );
  AND2X1_RVT U508 ( .A1(n26), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U509 ( .A1(n26), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U510 ( .A1(n26), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U511 ( .A1(n26), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U512 ( .A1(n26), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U513 ( .A1(n26), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U514 ( .A1(n26), .A2(n57), .Y(ab_16__0_) );
  AND2X1_RVT U515 ( .A1(n25), .A2(n75), .Y(ab_15__9_) );
  AND2X1_RVT U516 ( .A1(n25), .A2(n73), .Y(ab_15__8_) );
  AND2X1_RVT U517 ( .A1(n25), .A2(n71), .Y(ab_15__7_) );
  AND2X1_RVT U518 ( .A1(n25), .A2(n69), .Y(ab_15__6_) );
  AND2X1_RVT U519 ( .A1(n25), .A2(n67), .Y(ab_15__5_) );
  AND2X1_RVT U520 ( .A1(n25), .A2(n65), .Y(ab_15__4_) );
  AND2X1_RVT U521 ( .A1(A[15]), .A2(n62), .Y(ab_15__3_) );
  AND2X1_RVT U522 ( .A1(n25), .A2(n60), .Y(ab_15__2_) );
  AND2X1_RVT U523 ( .A1(A[15]), .A2(n58), .Y(ab_15__1_) );
  AND2X1_RVT U524 ( .A1(n25), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U525 ( .A1(n25), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U526 ( .A1(n25), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U527 ( .A1(n25), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U528 ( .A1(n25), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U529 ( .A1(n25), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U530 ( .A1(n25), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U531 ( .A1(A[15]), .A2(n57), .Y(ab_15__0_) );
  AND2X1_RVT U532 ( .A1(n24), .A2(n75), .Y(ab_14__9_) );
  AND2X1_RVT U533 ( .A1(n24), .A2(n73), .Y(ab_14__8_) );
  AND2X1_RVT U534 ( .A1(n24), .A2(n71), .Y(ab_14__7_) );
  AND2X1_RVT U535 ( .A1(n24), .A2(n69), .Y(ab_14__6_) );
  AND2X1_RVT U536 ( .A1(n24), .A2(n67), .Y(ab_14__5_) );
  AND2X1_RVT U537 ( .A1(A[14]), .A2(n65), .Y(ab_14__4_) );
  AND2X1_RVT U538 ( .A1(n24), .A2(n62), .Y(ab_14__3_) );
  AND2X1_RVT U539 ( .A1(A[14]), .A2(n60), .Y(ab_14__2_) );
  AND2X1_RVT U540 ( .A1(n24), .A2(n58), .Y(ab_14__1_) );
  AND2X1_RVT U541 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U542 ( .A1(n24), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U543 ( .A1(n24), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U544 ( .A1(n24), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U545 ( .A1(n24), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U546 ( .A1(n24), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U547 ( .A1(n24), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U548 ( .A1(n24), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U549 ( .A1(A[14]), .A2(n57), .Y(ab_14__0_) );
  AND2X1_RVT U550 ( .A1(n23), .A2(n75), .Y(ab_13__9_) );
  AND2X1_RVT U551 ( .A1(n23), .A2(n73), .Y(ab_13__8_) );
  AND2X1_RVT U552 ( .A1(A[13]), .A2(n71), .Y(ab_13__7_) );
  AND2X1_RVT U553 ( .A1(n23), .A2(n69), .Y(ab_13__6_) );
  AND2X1_RVT U554 ( .A1(A[13]), .A2(n67), .Y(ab_13__5_) );
  AND2X1_RVT U555 ( .A1(n23), .A2(n65), .Y(ab_13__4_) );
  AND2X1_RVT U556 ( .A1(A[13]), .A2(n62), .Y(ab_13__3_) );
  AND2X1_RVT U557 ( .A1(n23), .A2(n60), .Y(ab_13__2_) );
  AND2X1_RVT U558 ( .A1(A[13]), .A2(n58), .Y(ab_13__1_) );
  AND2X1_RVT U559 ( .A1(n23), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U560 ( .A1(n23), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U561 ( .A1(n23), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U562 ( .A1(n23), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U563 ( .A1(n23), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U564 ( .A1(n23), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U565 ( .A1(n23), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U566 ( .A1(n23), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U567 ( .A1(n23), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U568 ( .A1(A[13]), .A2(n57), .Y(ab_13__0_) );
  AND2X1_RVT U569 ( .A1(n22), .A2(n75), .Y(ab_12__9_) );
  AND2X1_RVT U570 ( .A1(n22), .A2(n73), .Y(ab_12__8_) );
  AND2X1_RVT U571 ( .A1(n22), .A2(n71), .Y(ab_12__7_) );
  AND2X1_RVT U572 ( .A1(A[12]), .A2(n69), .Y(ab_12__6_) );
  AND2X1_RVT U573 ( .A1(n22), .A2(n67), .Y(ab_12__5_) );
  AND2X1_RVT U574 ( .A1(A[12]), .A2(n65), .Y(ab_12__4_) );
  AND2X1_RVT U575 ( .A1(n22), .A2(n62), .Y(ab_12__3_) );
  AND2X1_RVT U576 ( .A1(A[12]), .A2(n60), .Y(ab_12__2_) );
  AND2X1_RVT U577 ( .A1(n22), .A2(n59), .Y(ab_12__1_) );
  AND2X1_RVT U578 ( .A1(A[12]), .A2(n14), .Y(ab_12__19_) );
  AND2X1_RVT U579 ( .A1(n22), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U580 ( .A1(n22), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U581 ( .A1(n22), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U582 ( .A1(n22), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U583 ( .A1(n22), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U584 ( .A1(n22), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U585 ( .A1(n22), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U586 ( .A1(n22), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U587 ( .A1(n22), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U588 ( .A1(A[12]), .A2(n57), .Y(ab_12__0_) );
  AND2X1_RVT U589 ( .A1(n21), .A2(n75), .Y(ab_11__9_) );
  AND2X1_RVT U590 ( .A1(n21), .A2(n73), .Y(ab_11__8_) );
  AND2X1_RVT U591 ( .A1(A[11]), .A2(n71), .Y(ab_11__7_) );
  AND2X1_RVT U592 ( .A1(n21), .A2(n69), .Y(ab_11__6_) );
  AND2X1_RVT U593 ( .A1(A[11]), .A2(n67), .Y(ab_11__5_) );
  AND2X1_RVT U594 ( .A1(n21), .A2(n65), .Y(ab_11__4_) );
  AND2X1_RVT U595 ( .A1(A[11]), .A2(n62), .Y(ab_11__3_) );
  AND2X1_RVT U596 ( .A1(n21), .A2(n61), .Y(ab_11__2_) );
  AND2X1_RVT U597 ( .A1(A[11]), .A2(n15), .Y(ab_11__20_) );
  AND2X1_RVT U598 ( .A1(n21), .A2(n59), .Y(ab_11__1_) );
  AND2X1_RVT U599 ( .A1(A[11]), .A2(n14), .Y(ab_11__19_) );
  AND2X1_RVT U600 ( .A1(n21), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U601 ( .A1(n21), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U602 ( .A1(n21), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U603 ( .A1(n21), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U604 ( .A1(n21), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U605 ( .A1(n21), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U606 ( .A1(n21), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U607 ( .A1(n21), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U608 ( .A1(n21), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U609 ( .A1(A[11]), .A2(n57), .Y(ab_11__0_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n75), .Y(ab_10__9_) );
  AND2X1_RVT U611 ( .A1(n20), .A2(n73), .Y(ab_10__8_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n71), .Y(ab_10__7_) );
  AND2X1_RVT U613 ( .A1(n20), .A2(n69), .Y(ab_10__6_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n67), .Y(ab_10__5_) );
  AND2X1_RVT U615 ( .A1(n20), .A2(n65), .Y(ab_10__4_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n63), .Y(ab_10__3_) );
  AND2X1_RVT U617 ( .A1(n20), .A2(n61), .Y(ab_10__2_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n16), .Y(ab_10__21_) );
  AND2X1_RVT U619 ( .A1(n20), .A2(n15), .Y(ab_10__20_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n59), .Y(ab_10__1_) );
  AND2X1_RVT U621 ( .A1(n20), .A2(n14), .Y(ab_10__19_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U623 ( .A1(n20), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U625 ( .A1(n20), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U627 ( .A1(n20), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U629 ( .A1(n20), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U631 ( .A1(n20), .A2(n57), .Y(ab_10__0_) );
  AND2X1_RVT U632 ( .A1(n36), .A2(n75), .Y(ab_0__9_) );
  AND2X1_RVT U633 ( .A1(n36), .A2(n73), .Y(ab_0__8_) );
  AND2X1_RVT U634 ( .A1(n36), .A2(n71), .Y(ab_0__7_) );
  AND2X1_RVT U635 ( .A1(n36), .A2(n69), .Y(ab_0__6_) );
  AND2X1_RVT U636 ( .A1(n36), .A2(n67), .Y(ab_0__5_) );
  AND2X1_RVT U637 ( .A1(n36), .A2(n64), .Y(ab_0__4_) );
  AND2X1_RVT U638 ( .A1(n36), .A2(n63), .Y(ab_0__3_) );
  AND2X1_RVT U639 ( .A1(n36), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U640 ( .A1(n35), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U641 ( .A1(n35), .A2(n61), .Y(ab_0__2_) );
  AND2X1_RVT U642 ( .A1(n35), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U643 ( .A1(n35), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U644 ( .A1(n35), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U645 ( .A1(n35), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U646 ( .A1(n35), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U647 ( .A1(n35), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U648 ( .A1(n35), .A2(n18), .Y(ab_0__23_) );
  AND2X1_RVT U649 ( .A1(n35), .A2(n17), .Y(ab_0__22_) );
  AND2X1_RVT U650 ( .A1(n35), .A2(n16), .Y(ab_0__21_) );
  AND2X1_RVT U651 ( .A1(n35), .A2(n15), .Y(ab_0__20_) );
  AND2X1_RVT U652 ( .A1(n34), .A2(n59), .Y(ab_0__1_) );
  AND2X1_RVT U653 ( .A1(n34), .A2(n14), .Y(ab_0__19_) );
  AND2X1_RVT U654 ( .A1(n34), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U655 ( .A1(n34), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U656 ( .A1(n34), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U657 ( .A1(n34), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U658 ( .A1(n34), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U659 ( .A1(n34), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U660 ( .A1(n34), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U661 ( .A1(n34), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U662 ( .A1(n34), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U663 ( .A1(n34), .A2(n57), .Y(PRODUCT_0_) );
endmodule


module OSPE_14_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_14 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n2), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n3), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n4), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n4), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n4), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n4), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n4), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n4), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n2), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n3), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n4), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n1), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n1), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n1), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n1), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n1), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n1), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n1), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n1), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n1), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n1), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n1), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n1), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n1), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n1), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n2), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n2), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n2), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n2), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n2), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n2), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n2), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n2), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n2), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n2), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n2), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n2), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_14_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_14_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_13_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U5 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U6 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U7 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U8 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U9 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U10 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U11 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U12 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U13 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U14 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U15 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U16 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U17 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U18 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U19 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U20 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U21 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  XOR2X1_RVT U22 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U23 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U24 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR2X1_RVT U25 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U27 ( .A(A[1]), .Y(n38) );
  NBUFFX2_RVT U28 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U29 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U30 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U31 ( .A(A[3]), .Y(n42) );
  XOR2X1_RVT U32 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U33 ( .A(A[0]), .Y(n36) );
  NBUFFX2_RVT U34 ( .A(A[1]), .Y(n39) );
  XOR2X1_RVT U35 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U36 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U37 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U38 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U39 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n41) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n63) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n75) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n73) );
  NBUFFX2_RVT U44 ( .A(B[7]), .Y(n71) );
  NBUFFX2_RVT U45 ( .A(A[9]), .Y(n55) );
  NBUFFX2_RVT U46 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U47 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U48 ( .A(B[6]), .Y(n69) );
  NBUFFX2_RVT U49 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U50 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U51 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U52 ( .A(B[5]), .Y(n66) );
  NBUFFX2_RVT U53 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U54 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U55 ( .A(B[4]), .Y(n65) );
  NBUFFX2_RVT U56 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U57 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U58 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U59 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U60 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U61 ( .A(A[6]), .Y(n48) );
  NBUFFX2_RVT U62 ( .A(A[7]), .Y(n51) );
  NBUFFX2_RVT U63 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U64 ( .A(B[5]), .Y(n67) );
  NBUFFX2_RVT U65 ( .A(A[8]), .Y(n53) );
  NBUFFX2_RVT U66 ( .A(A[8]), .Y(n52) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n43) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n57) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n45) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n59) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n47) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n61) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n49) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  NBUFFX2_RVT U116 ( .A(B[19]), .Y(n14) );
  NBUFFX2_RVT U117 ( .A(B[20]), .Y(n15) );
  NBUFFX2_RVT U118 ( .A(B[21]), .Y(n16) );
  NBUFFX2_RVT U119 ( .A(B[22]), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(B[23]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[10]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[11]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[12]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[13]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[14]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[15]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[16]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[17]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[18]), .Y(n28) );
  NBUFFX2_RVT U131 ( .A(A[19]), .Y(n29) );
  INVX0_RVT U132 ( .A(A[20]), .Y(n30) );
  INVX0_RVT U133 ( .A(n30), .Y(n31) );
  INVX0_RVT U134 ( .A(A[21]), .Y(n32) );
  INVX0_RVT U135 ( .A(n32), .Y(n33) );
  AND2X1_RVT U136 ( .A1(n74), .A2(n55), .Y(ab_9__9_) );
  AND2X1_RVT U137 ( .A1(n72), .A2(n55), .Y(ab_9__8_) );
  AND2X1_RVT U138 ( .A1(n70), .A2(n55), .Y(ab_9__7_) );
  AND2X1_RVT U139 ( .A1(n68), .A2(n55), .Y(ab_9__6_) );
  AND2X1_RVT U140 ( .A1(n66), .A2(n55), .Y(ab_9__5_) );
  AND2X1_RVT U141 ( .A1(n64), .A2(n55), .Y(ab_9__4_) );
  AND2X1_RVT U142 ( .A1(n63), .A2(n55), .Y(ab_9__3_) );
  AND2X1_RVT U143 ( .A1(n61), .A2(n55), .Y(ab_9__2_) );
  AND2X1_RVT U144 ( .A1(n17), .A2(n55), .Y(ab_9__22_) );
  AND2X1_RVT U145 ( .A1(n16), .A2(n55), .Y(ab_9__21_) );
  AND2X1_RVT U146 ( .A1(n15), .A2(n55), .Y(ab_9__20_) );
  AND2X1_RVT U147 ( .A1(n59), .A2(n54), .Y(ab_9__1_) );
  AND2X1_RVT U148 ( .A1(n14), .A2(n54), .Y(ab_9__19_) );
  AND2X1_RVT U149 ( .A1(n13), .A2(n54), .Y(ab_9__18_) );
  AND2X1_RVT U150 ( .A1(B[17]), .A2(n54), .Y(ab_9__17_) );
  AND2X1_RVT U151 ( .A1(n11), .A2(n54), .Y(ab_9__16_) );
  AND2X1_RVT U152 ( .A1(n10), .A2(n54), .Y(ab_9__15_) );
  AND2X1_RVT U153 ( .A1(n9), .A2(n54), .Y(ab_9__14_) );
  AND2X1_RVT U154 ( .A1(B[13]), .A2(n54), .Y(ab_9__13_) );
  AND2X1_RVT U155 ( .A1(n7), .A2(n54), .Y(ab_9__12_) );
  AND2X1_RVT U156 ( .A1(n5), .A2(n54), .Y(ab_9__11_) );
  AND2X1_RVT U157 ( .A1(n3), .A2(n54), .Y(ab_9__10_) );
  AND2X1_RVT U158 ( .A1(n56), .A2(n54), .Y(ab_9__0_) );
  AND2X1_RVT U159 ( .A1(n53), .A2(n74), .Y(ab_8__9_) );
  AND2X1_RVT U160 ( .A1(n53), .A2(n72), .Y(ab_8__8_) );
  AND2X1_RVT U161 ( .A1(n53), .A2(n70), .Y(ab_8__7_) );
  AND2X1_RVT U162 ( .A1(n53), .A2(n68), .Y(ab_8__6_) );
  AND2X1_RVT U163 ( .A1(n53), .A2(n66), .Y(ab_8__5_) );
  AND2X1_RVT U164 ( .A1(n53), .A2(n64), .Y(ab_8__4_) );
  AND2X1_RVT U165 ( .A1(n53), .A2(n63), .Y(ab_8__3_) );
  AND2X1_RVT U166 ( .A1(n53), .A2(n61), .Y(ab_8__2_) );
  AND2X1_RVT U167 ( .A1(n53), .A2(n18), .Y(ab_8__23_) );
  AND2X1_RVT U168 ( .A1(n53), .A2(n17), .Y(ab_8__22_) );
  AND2X1_RVT U169 ( .A1(n53), .A2(n16), .Y(ab_8__21_) );
  AND2X1_RVT U170 ( .A1(n53), .A2(n15), .Y(ab_8__20_) );
  AND2X1_RVT U171 ( .A1(n52), .A2(n59), .Y(ab_8__1_) );
  AND2X1_RVT U172 ( .A1(n52), .A2(n14), .Y(ab_8__19_) );
  AND2X1_RVT U173 ( .A1(n52), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U174 ( .A1(n52), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U175 ( .A1(n52), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U176 ( .A1(n52), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U177 ( .A1(n52), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U178 ( .A1(n52), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U179 ( .A1(n52), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U180 ( .A1(n52), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U181 ( .A1(n52), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U182 ( .A1(n52), .A2(n56), .Y(ab_8__0_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n74), .Y(ab_7__9_) );
  AND2X1_RVT U184 ( .A1(n51), .A2(n72), .Y(ab_7__8_) );
  AND2X1_RVT U185 ( .A1(n51), .A2(n70), .Y(ab_7__7_) );
  AND2X1_RVT U186 ( .A1(n51), .A2(n68), .Y(ab_7__6_) );
  AND2X1_RVT U187 ( .A1(n51), .A2(n66), .Y(ab_7__5_) );
  AND2X1_RVT U188 ( .A1(n51), .A2(n64), .Y(ab_7__4_) );
  AND2X1_RVT U189 ( .A1(n51), .A2(n63), .Y(ab_7__3_) );
  AND2X1_RVT U190 ( .A1(n51), .A2(n61), .Y(ab_7__2_) );
  AND2X1_RVT U191 ( .A1(n51), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U192 ( .A1(n51), .A2(n18), .Y(ab_7__23_) );
  AND2X1_RVT U193 ( .A1(n51), .A2(n17), .Y(ab_7__22_) );
  AND2X1_RVT U194 ( .A1(n51), .A2(n16), .Y(ab_7__21_) );
  AND2X1_RVT U195 ( .A1(n51), .A2(n15), .Y(ab_7__20_) );
  AND2X1_RVT U196 ( .A1(n50), .A2(n59), .Y(ab_7__1_) );
  AND2X1_RVT U197 ( .A1(n50), .A2(n14), .Y(ab_7__19_) );
  AND2X1_RVT U198 ( .A1(n50), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U199 ( .A1(n50), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U200 ( .A1(n50), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U201 ( .A1(n50), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U202 ( .A1(n50), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U203 ( .A1(n50), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U204 ( .A1(n50), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U205 ( .A1(n50), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U206 ( .A1(n50), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U207 ( .A1(n50), .A2(n56), .Y(ab_7__0_) );
  AND2X1_RVT U208 ( .A1(n49), .A2(n74), .Y(ab_6__9_) );
  AND2X1_RVT U209 ( .A1(n49), .A2(n72), .Y(ab_6__8_) );
  AND2X1_RVT U210 ( .A1(n48), .A2(n70), .Y(ab_6__7_) );
  AND2X1_RVT U211 ( .A1(n48), .A2(n68), .Y(ab_6__6_) );
  AND2X1_RVT U212 ( .A1(n48), .A2(n66), .Y(ab_6__5_) );
  AND2X1_RVT U213 ( .A1(n48), .A2(n64), .Y(ab_6__4_) );
  AND2X1_RVT U214 ( .A1(n48), .A2(n63), .Y(ab_6__3_) );
  AND2X1_RVT U215 ( .A1(n48), .A2(n61), .Y(ab_6__2_) );
  AND2X1_RVT U216 ( .A1(n48), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U217 ( .A1(n48), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U218 ( .A1(n48), .A2(n18), .Y(ab_6__23_) );
  AND2X1_RVT U219 ( .A1(n48), .A2(n17), .Y(ab_6__22_) );
  AND2X1_RVT U220 ( .A1(n48), .A2(n16), .Y(ab_6__21_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n15), .Y(ab_6__20_) );
  AND2X1_RVT U222 ( .A1(n49), .A2(n59), .Y(ab_6__1_) );
  AND2X1_RVT U223 ( .A1(n49), .A2(n14), .Y(ab_6__19_) );
  AND2X1_RVT U224 ( .A1(n49), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U225 ( .A1(n49), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U226 ( .A1(n49), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U227 ( .A1(n49), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U228 ( .A1(n49), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U229 ( .A1(n49), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U230 ( .A1(n49), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U231 ( .A1(n49), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U232 ( .A1(n49), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U233 ( .A1(n49), .A2(n56), .Y(ab_6__0_) );
  AND2X1_RVT U234 ( .A1(n47), .A2(n74), .Y(ab_5__9_) );
  AND2X1_RVT U235 ( .A1(n47), .A2(n72), .Y(ab_5__8_) );
  AND2X1_RVT U236 ( .A1(n47), .A2(n70), .Y(ab_5__7_) );
  AND2X1_RVT U237 ( .A1(n46), .A2(n68), .Y(ab_5__6_) );
  AND2X1_RVT U238 ( .A1(n46), .A2(n66), .Y(ab_5__5_) );
  AND2X1_RVT U239 ( .A1(n46), .A2(n64), .Y(ab_5__4_) );
  AND2X1_RVT U240 ( .A1(n46), .A2(n63), .Y(ab_5__3_) );
  AND2X1_RVT U241 ( .A1(n46), .A2(n61), .Y(ab_5__2_) );
  AND2X1_RVT U242 ( .A1(n46), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U243 ( .A1(n46), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U244 ( .A1(n46), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U245 ( .A1(n46), .A2(n18), .Y(ab_5__23_) );
  AND2X1_RVT U246 ( .A1(n46), .A2(n17), .Y(ab_5__22_) );
  AND2X1_RVT U247 ( .A1(n46), .A2(n16), .Y(ab_5__21_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n15), .Y(ab_5__20_) );
  AND2X1_RVT U249 ( .A1(n47), .A2(n59), .Y(ab_5__1_) );
  AND2X1_RVT U250 ( .A1(n47), .A2(n14), .Y(ab_5__19_) );
  AND2X1_RVT U251 ( .A1(n47), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U252 ( .A1(n47), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U253 ( .A1(n47), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U254 ( .A1(n47), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U255 ( .A1(n47), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U256 ( .A1(n47), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U257 ( .A1(n47), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U258 ( .A1(n47), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U259 ( .A1(n47), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U260 ( .A1(n47), .A2(n56), .Y(ab_5__0_) );
  AND2X1_RVT U261 ( .A1(n45), .A2(n74), .Y(ab_4__9_) );
  AND2X1_RVT U262 ( .A1(n45), .A2(n72), .Y(ab_4__8_) );
  AND2X1_RVT U263 ( .A1(n45), .A2(n70), .Y(ab_4__7_) );
  AND2X1_RVT U264 ( .A1(n45), .A2(n68), .Y(ab_4__6_) );
  AND2X1_RVT U265 ( .A1(n44), .A2(n66), .Y(ab_4__5_) );
  AND2X1_RVT U266 ( .A1(n44), .A2(n64), .Y(ab_4__4_) );
  AND2X1_RVT U267 ( .A1(n44), .A2(n63), .Y(ab_4__3_) );
  AND2X1_RVT U268 ( .A1(n44), .A2(n61), .Y(ab_4__2_) );
  AND2X1_RVT U269 ( .A1(n44), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U270 ( .A1(n44), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U271 ( .A1(n44), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U272 ( .A1(n44), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U273 ( .A1(n44), .A2(n18), .Y(ab_4__23_) );
  AND2X1_RVT U274 ( .A1(n44), .A2(n17), .Y(ab_4__22_) );
  AND2X1_RVT U275 ( .A1(n44), .A2(n16), .Y(ab_4__21_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n15), .Y(ab_4__20_) );
  AND2X1_RVT U277 ( .A1(n45), .A2(n59), .Y(ab_4__1_) );
  AND2X1_RVT U278 ( .A1(n45), .A2(n14), .Y(ab_4__19_) );
  AND2X1_RVT U279 ( .A1(n45), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U280 ( .A1(n45), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U281 ( .A1(n45), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U282 ( .A1(n45), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U283 ( .A1(n45), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U284 ( .A1(n45), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U285 ( .A1(n45), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U286 ( .A1(n45), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U287 ( .A1(n45), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U288 ( .A1(n45), .A2(n56), .Y(ab_4__0_) );
  AND2X1_RVT U289 ( .A1(n43), .A2(n74), .Y(ab_3__9_) );
  AND2X1_RVT U290 ( .A1(n43), .A2(n72), .Y(ab_3__8_) );
  AND2X1_RVT U291 ( .A1(n43), .A2(n70), .Y(ab_3__7_) );
  AND2X1_RVT U292 ( .A1(n43), .A2(n68), .Y(ab_3__6_) );
  AND2X1_RVT U293 ( .A1(n43), .A2(n66), .Y(ab_3__5_) );
  AND2X1_RVT U294 ( .A1(n42), .A2(n64), .Y(ab_3__4_) );
  AND2X1_RVT U295 ( .A1(n42), .A2(n63), .Y(ab_3__3_) );
  AND2X1_RVT U296 ( .A1(n42), .A2(n61), .Y(ab_3__2_) );
  AND2X1_RVT U297 ( .A1(n42), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U298 ( .A1(n42), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U299 ( .A1(n42), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U300 ( .A1(n42), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U301 ( .A1(n42), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U302 ( .A1(n42), .A2(n18), .Y(ab_3__23_) );
  AND2X1_RVT U303 ( .A1(n42), .A2(n17), .Y(ab_3__22_) );
  AND2X1_RVT U304 ( .A1(n42), .A2(n16), .Y(ab_3__21_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n15), .Y(ab_3__20_) );
  AND2X1_RVT U306 ( .A1(n43), .A2(n59), .Y(ab_3__1_) );
  AND2X1_RVT U307 ( .A1(n43), .A2(n14), .Y(ab_3__19_) );
  AND2X1_RVT U308 ( .A1(n43), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U309 ( .A1(n43), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U310 ( .A1(n43), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U311 ( .A1(n43), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U312 ( .A1(n43), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U313 ( .A1(n43), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U314 ( .A1(n43), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U315 ( .A1(n43), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U316 ( .A1(n43), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U317 ( .A1(n43), .A2(n56), .Y(ab_3__0_) );
  AND2X1_RVT U318 ( .A1(A[31]), .A2(n56), .Y(ab_31__0_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n59), .Y(ab_30__1_) );
  AND2X1_RVT U320 ( .A1(A[30]), .A2(n56), .Y(ab_30__0_) );
  AND2X1_RVT U321 ( .A1(n41), .A2(n74), .Y(ab_2__9_) );
  AND2X1_RVT U322 ( .A1(n41), .A2(n72), .Y(ab_2__8_) );
  AND2X1_RVT U323 ( .A1(n41), .A2(n70), .Y(ab_2__7_) );
  AND2X1_RVT U324 ( .A1(n41), .A2(n68), .Y(ab_2__6_) );
  AND2X1_RVT U325 ( .A1(n41), .A2(n66), .Y(ab_2__5_) );
  AND2X1_RVT U326 ( .A1(n41), .A2(n64), .Y(ab_2__4_) );
  AND2X1_RVT U327 ( .A1(n41), .A2(n63), .Y(ab_2__3_) );
  AND2X1_RVT U328 ( .A1(n40), .A2(n61), .Y(ab_2__2_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U330 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U331 ( .A1(n41), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U332 ( .A1(n40), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U333 ( .A1(n40), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U334 ( .A1(n40), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U335 ( .A1(A[2]), .A2(n18), .Y(ab_2__23_) );
  AND2X1_RVT U336 ( .A1(n41), .A2(n17), .Y(ab_2__22_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n16), .Y(ab_2__21_) );
  AND2X1_RVT U338 ( .A1(A[2]), .A2(n15), .Y(ab_2__20_) );
  AND2X1_RVT U339 ( .A1(n40), .A2(n59), .Y(ab_2__1_) );
  AND2X1_RVT U340 ( .A1(n40), .A2(n14), .Y(ab_2__19_) );
  AND2X1_RVT U341 ( .A1(n40), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U342 ( .A1(n40), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U343 ( .A1(n40), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U344 ( .A1(n40), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U345 ( .A1(n40), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U346 ( .A1(n40), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U347 ( .A1(n40), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U348 ( .A1(n40), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U349 ( .A1(n40), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U350 ( .A1(n40), .A2(n56), .Y(ab_2__0_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n61), .Y(ab_29__2_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n59), .Y(ab_29__1_) );
  AND2X1_RVT U353 ( .A1(A[29]), .A2(n56), .Y(ab_29__0_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n63), .Y(ab_28__3_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n61), .Y(ab_28__2_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n59), .Y(ab_28__1_) );
  AND2X1_RVT U357 ( .A1(A[28]), .A2(n56), .Y(ab_28__0_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n64), .Y(ab_27__4_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n63), .Y(ab_27__3_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n61), .Y(ab_27__2_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n59), .Y(ab_27__1_) );
  AND2X1_RVT U362 ( .A1(A[27]), .A2(n56), .Y(ab_27__0_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n66), .Y(ab_26__5_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n64), .Y(ab_26__4_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n63), .Y(ab_26__3_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n61), .Y(ab_26__2_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n59), .Y(ab_26__1_) );
  AND2X1_RVT U368 ( .A1(A[26]), .A2(n57), .Y(ab_26__0_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n68), .Y(ab_25__6_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n66), .Y(ab_25__5_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n64), .Y(ab_25__4_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n63), .Y(ab_25__3_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n61), .Y(ab_25__2_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n58), .Y(ab_25__1_) );
  AND2X1_RVT U375 ( .A1(A[25]), .A2(n57), .Y(ab_25__0_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n70), .Y(ab_24__7_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n68), .Y(ab_24__6_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n66), .Y(ab_24__5_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n64), .Y(ab_24__4_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n63), .Y(ab_24__3_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n60), .Y(ab_24__2_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n58), .Y(ab_24__1_) );
  AND2X1_RVT U383 ( .A1(A[24]), .A2(n57), .Y(ab_24__0_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n72), .Y(ab_23__8_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n70), .Y(ab_23__7_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n68), .Y(ab_23__6_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n66), .Y(ab_23__5_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n64), .Y(ab_23__4_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n62), .Y(ab_23__3_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n60), .Y(ab_23__2_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n58), .Y(ab_23__1_) );
  AND2X1_RVT U392 ( .A1(A[23]), .A2(n57), .Y(ab_23__0_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n74), .Y(ab_22__9_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n72), .Y(ab_22__8_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n70), .Y(ab_22__7_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n68), .Y(ab_22__6_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n66), .Y(ab_22__5_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n65), .Y(ab_22__4_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n62), .Y(ab_22__3_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n60), .Y(ab_22__2_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n58), .Y(ab_22__1_) );
  AND2X1_RVT U402 ( .A1(A[22]), .A2(n57), .Y(ab_22__0_) );
  AND2X1_RVT U403 ( .A1(A[21]), .A2(n74), .Y(ab_21__9_) );
  AND2X1_RVT U404 ( .A1(n33), .A2(n72), .Y(ab_21__8_) );
  AND2X1_RVT U405 ( .A1(n33), .A2(n70), .Y(ab_21__7_) );
  AND2X1_RVT U406 ( .A1(n33), .A2(n68), .Y(ab_21__6_) );
  AND2X1_RVT U407 ( .A1(n33), .A2(n67), .Y(ab_21__5_) );
  AND2X1_RVT U408 ( .A1(n33), .A2(n65), .Y(ab_21__4_) );
  AND2X1_RVT U409 ( .A1(n33), .A2(n62), .Y(ab_21__3_) );
  AND2X1_RVT U410 ( .A1(n33), .A2(n60), .Y(ab_21__2_) );
  AND2X1_RVT U411 ( .A1(n33), .A2(n58), .Y(ab_21__1_) );
  AND2X1_RVT U412 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U413 ( .A1(n33), .A2(n57), .Y(ab_21__0_) );
  AND2X1_RVT U414 ( .A1(n31), .A2(n74), .Y(ab_20__9_) );
  AND2X1_RVT U415 ( .A1(n31), .A2(n72), .Y(ab_20__8_) );
  AND2X1_RVT U416 ( .A1(n31), .A2(n70), .Y(ab_20__7_) );
  AND2X1_RVT U417 ( .A1(n31), .A2(n69), .Y(ab_20__6_) );
  AND2X1_RVT U418 ( .A1(n31), .A2(n67), .Y(ab_20__5_) );
  AND2X1_RVT U419 ( .A1(n31), .A2(n65), .Y(ab_20__4_) );
  AND2X1_RVT U420 ( .A1(n31), .A2(n62), .Y(ab_20__3_) );
  AND2X1_RVT U421 ( .A1(n31), .A2(n60), .Y(ab_20__2_) );
  AND2X1_RVT U422 ( .A1(n31), .A2(n58), .Y(ab_20__1_) );
  AND2X1_RVT U423 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U424 ( .A1(n31), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U425 ( .A1(n31), .A2(n57), .Y(ab_20__0_) );
  AND2X1_RVT U426 ( .A1(n39), .A2(n74), .Y(ab_1__9_) );
  AND2X1_RVT U427 ( .A1(n39), .A2(n72), .Y(ab_1__8_) );
  AND2X1_RVT U428 ( .A1(n39), .A2(n71), .Y(ab_1__7_) );
  AND2X1_RVT U429 ( .A1(n39), .A2(n69), .Y(ab_1__6_) );
  AND2X1_RVT U430 ( .A1(n39), .A2(n67), .Y(ab_1__5_) );
  AND2X1_RVT U431 ( .A1(n39), .A2(n65), .Y(ab_1__4_) );
  AND2X1_RVT U432 ( .A1(n39), .A2(n62), .Y(ab_1__3_) );
  AND2X1_RVT U433 ( .A1(n38), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U434 ( .A1(n38), .A2(n60), .Y(ab_1__2_) );
  AND2X1_RVT U435 ( .A1(n38), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U436 ( .A1(n38), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U437 ( .A1(n38), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U438 ( .A1(n38), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U439 ( .A1(n38), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U440 ( .A1(n38), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U441 ( .A1(n38), .A2(n18), .Y(ab_1__23_) );
  AND2X1_RVT U442 ( .A1(n38), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U443 ( .A1(n38), .A2(n16), .Y(ab_1__21_) );
  AND2X1_RVT U444 ( .A1(n38), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U445 ( .A1(n37), .A2(n58), .Y(ab_1__1_) );
  AND2X1_RVT U446 ( .A1(n37), .A2(n14), .Y(ab_1__19_) );
  AND2X1_RVT U447 ( .A1(n37), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U448 ( .A1(n37), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U449 ( .A1(n37), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U450 ( .A1(n37), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U451 ( .A1(n37), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U452 ( .A1(n37), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U453 ( .A1(n37), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U454 ( .A1(n37), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U455 ( .A1(n37), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U456 ( .A1(n37), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U457 ( .A1(n29), .A2(n74), .Y(ab_19__9_) );
  AND2X1_RVT U458 ( .A1(n29), .A2(n73), .Y(ab_19__8_) );
  AND2X1_RVT U459 ( .A1(n29), .A2(n71), .Y(ab_19__7_) );
  AND2X1_RVT U460 ( .A1(n29), .A2(n69), .Y(ab_19__6_) );
  AND2X1_RVT U461 ( .A1(n29), .A2(n67), .Y(ab_19__5_) );
  AND2X1_RVT U462 ( .A1(n29), .A2(n65), .Y(ab_19__4_) );
  AND2X1_RVT U463 ( .A1(n29), .A2(n62), .Y(ab_19__3_) );
  AND2X1_RVT U464 ( .A1(n29), .A2(n60), .Y(ab_19__2_) );
  AND2X1_RVT U465 ( .A1(n29), .A2(n58), .Y(ab_19__1_) );
  AND2X1_RVT U466 ( .A1(n29), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U467 ( .A1(n29), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U468 ( .A1(n29), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U469 ( .A1(A[19]), .A2(n57), .Y(ab_19__0_) );
  AND2X1_RVT U470 ( .A1(n28), .A2(n75), .Y(ab_18__9_) );
  AND2X1_RVT U471 ( .A1(n28), .A2(n73), .Y(ab_18__8_) );
  AND2X1_RVT U472 ( .A1(n28), .A2(n71), .Y(ab_18__7_) );
  AND2X1_RVT U473 ( .A1(n28), .A2(n69), .Y(ab_18__6_) );
  AND2X1_RVT U474 ( .A1(n28), .A2(n67), .Y(ab_18__5_) );
  AND2X1_RVT U475 ( .A1(n28), .A2(n65), .Y(ab_18__4_) );
  AND2X1_RVT U476 ( .A1(n28), .A2(n62), .Y(ab_18__3_) );
  AND2X1_RVT U477 ( .A1(n28), .A2(n60), .Y(ab_18__2_) );
  AND2X1_RVT U478 ( .A1(n28), .A2(n58), .Y(ab_18__1_) );
  AND2X1_RVT U479 ( .A1(A[18]), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U480 ( .A1(n28), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U481 ( .A1(n28), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U482 ( .A1(n28), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U483 ( .A1(n28), .A2(n57), .Y(ab_18__0_) );
  AND2X1_RVT U484 ( .A1(n27), .A2(n75), .Y(ab_17__9_) );
  AND2X1_RVT U485 ( .A1(n27), .A2(n73), .Y(ab_17__8_) );
  AND2X1_RVT U486 ( .A1(n27), .A2(n71), .Y(ab_17__7_) );
  AND2X1_RVT U487 ( .A1(n27), .A2(n69), .Y(ab_17__6_) );
  AND2X1_RVT U488 ( .A1(n27), .A2(n67), .Y(ab_17__5_) );
  AND2X1_RVT U489 ( .A1(n27), .A2(n65), .Y(ab_17__4_) );
  AND2X1_RVT U490 ( .A1(n27), .A2(n62), .Y(ab_17__3_) );
  AND2X1_RVT U491 ( .A1(n27), .A2(n60), .Y(ab_17__2_) );
  AND2X1_RVT U492 ( .A1(A[17]), .A2(n58), .Y(ab_17__1_) );
  AND2X1_RVT U493 ( .A1(n27), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U494 ( .A1(n27), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U495 ( .A1(n27), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U496 ( .A1(n27), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U497 ( .A1(n27), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U498 ( .A1(A[17]), .A2(n57), .Y(ab_17__0_) );
  AND2X1_RVT U499 ( .A1(n26), .A2(n75), .Y(ab_16__9_) );
  AND2X1_RVT U500 ( .A1(n26), .A2(n73), .Y(ab_16__8_) );
  AND2X1_RVT U501 ( .A1(n26), .A2(n71), .Y(ab_16__7_) );
  AND2X1_RVT U502 ( .A1(n26), .A2(n69), .Y(ab_16__6_) );
  AND2X1_RVT U503 ( .A1(n26), .A2(n67), .Y(ab_16__5_) );
  AND2X1_RVT U504 ( .A1(n26), .A2(n65), .Y(ab_16__4_) );
  AND2X1_RVT U505 ( .A1(A[16]), .A2(n62), .Y(ab_16__3_) );
  AND2X1_RVT U506 ( .A1(n26), .A2(n60), .Y(ab_16__2_) );
  AND2X1_RVT U507 ( .A1(A[16]), .A2(n58), .Y(ab_16__1_) );
  AND2X1_RVT U508 ( .A1(n26), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U509 ( .A1(n26), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U510 ( .A1(n26), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U511 ( .A1(n26), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U512 ( .A1(n26), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U513 ( .A1(n26), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U514 ( .A1(n26), .A2(n57), .Y(ab_16__0_) );
  AND2X1_RVT U515 ( .A1(n25), .A2(n75), .Y(ab_15__9_) );
  AND2X1_RVT U516 ( .A1(n25), .A2(n73), .Y(ab_15__8_) );
  AND2X1_RVT U517 ( .A1(n25), .A2(n71), .Y(ab_15__7_) );
  AND2X1_RVT U518 ( .A1(n25), .A2(n69), .Y(ab_15__6_) );
  AND2X1_RVT U519 ( .A1(n25), .A2(n67), .Y(ab_15__5_) );
  AND2X1_RVT U520 ( .A1(n25), .A2(n65), .Y(ab_15__4_) );
  AND2X1_RVT U521 ( .A1(A[15]), .A2(n62), .Y(ab_15__3_) );
  AND2X1_RVT U522 ( .A1(n25), .A2(n60), .Y(ab_15__2_) );
  AND2X1_RVT U523 ( .A1(A[15]), .A2(n58), .Y(ab_15__1_) );
  AND2X1_RVT U524 ( .A1(n25), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U525 ( .A1(n25), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U526 ( .A1(n25), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U527 ( .A1(n25), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U528 ( .A1(n25), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U529 ( .A1(n25), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U530 ( .A1(n25), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U531 ( .A1(A[15]), .A2(n57), .Y(ab_15__0_) );
  AND2X1_RVT U532 ( .A1(n24), .A2(n75), .Y(ab_14__9_) );
  AND2X1_RVT U533 ( .A1(n24), .A2(n73), .Y(ab_14__8_) );
  AND2X1_RVT U534 ( .A1(n24), .A2(n71), .Y(ab_14__7_) );
  AND2X1_RVT U535 ( .A1(n24), .A2(n69), .Y(ab_14__6_) );
  AND2X1_RVT U536 ( .A1(n24), .A2(n67), .Y(ab_14__5_) );
  AND2X1_RVT U537 ( .A1(A[14]), .A2(n65), .Y(ab_14__4_) );
  AND2X1_RVT U538 ( .A1(n24), .A2(n62), .Y(ab_14__3_) );
  AND2X1_RVT U539 ( .A1(A[14]), .A2(n60), .Y(ab_14__2_) );
  AND2X1_RVT U540 ( .A1(n24), .A2(n58), .Y(ab_14__1_) );
  AND2X1_RVT U541 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U542 ( .A1(n24), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U543 ( .A1(n24), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U544 ( .A1(n24), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U545 ( .A1(n24), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U546 ( .A1(n24), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U547 ( .A1(n24), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U548 ( .A1(n24), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U549 ( .A1(A[14]), .A2(n57), .Y(ab_14__0_) );
  AND2X1_RVT U550 ( .A1(n23), .A2(n75), .Y(ab_13__9_) );
  AND2X1_RVT U551 ( .A1(n23), .A2(n73), .Y(ab_13__8_) );
  AND2X1_RVT U552 ( .A1(A[13]), .A2(n71), .Y(ab_13__7_) );
  AND2X1_RVT U553 ( .A1(n23), .A2(n69), .Y(ab_13__6_) );
  AND2X1_RVT U554 ( .A1(A[13]), .A2(n67), .Y(ab_13__5_) );
  AND2X1_RVT U555 ( .A1(n23), .A2(n65), .Y(ab_13__4_) );
  AND2X1_RVT U556 ( .A1(A[13]), .A2(n62), .Y(ab_13__3_) );
  AND2X1_RVT U557 ( .A1(n23), .A2(n60), .Y(ab_13__2_) );
  AND2X1_RVT U558 ( .A1(A[13]), .A2(n58), .Y(ab_13__1_) );
  AND2X1_RVT U559 ( .A1(n23), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U560 ( .A1(n23), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U561 ( .A1(n23), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U562 ( .A1(n23), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U563 ( .A1(n23), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U564 ( .A1(n23), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U565 ( .A1(n23), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U566 ( .A1(n23), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U567 ( .A1(n23), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U568 ( .A1(A[13]), .A2(n57), .Y(ab_13__0_) );
  AND2X1_RVT U569 ( .A1(n22), .A2(n75), .Y(ab_12__9_) );
  AND2X1_RVT U570 ( .A1(n22), .A2(n73), .Y(ab_12__8_) );
  AND2X1_RVT U571 ( .A1(n22), .A2(n71), .Y(ab_12__7_) );
  AND2X1_RVT U572 ( .A1(A[12]), .A2(n69), .Y(ab_12__6_) );
  AND2X1_RVT U573 ( .A1(n22), .A2(n67), .Y(ab_12__5_) );
  AND2X1_RVT U574 ( .A1(A[12]), .A2(n65), .Y(ab_12__4_) );
  AND2X1_RVT U575 ( .A1(n22), .A2(n62), .Y(ab_12__3_) );
  AND2X1_RVT U576 ( .A1(A[12]), .A2(n60), .Y(ab_12__2_) );
  AND2X1_RVT U577 ( .A1(n22), .A2(n59), .Y(ab_12__1_) );
  AND2X1_RVT U578 ( .A1(A[12]), .A2(n14), .Y(ab_12__19_) );
  AND2X1_RVT U579 ( .A1(n22), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U580 ( .A1(n22), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U581 ( .A1(n22), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U582 ( .A1(n22), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U583 ( .A1(n22), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U584 ( .A1(n22), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U585 ( .A1(n22), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U586 ( .A1(n22), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U587 ( .A1(n22), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U588 ( .A1(A[12]), .A2(n57), .Y(ab_12__0_) );
  AND2X1_RVT U589 ( .A1(n21), .A2(n75), .Y(ab_11__9_) );
  AND2X1_RVT U590 ( .A1(n21), .A2(n73), .Y(ab_11__8_) );
  AND2X1_RVT U591 ( .A1(A[11]), .A2(n71), .Y(ab_11__7_) );
  AND2X1_RVT U592 ( .A1(n21), .A2(n69), .Y(ab_11__6_) );
  AND2X1_RVT U593 ( .A1(A[11]), .A2(n67), .Y(ab_11__5_) );
  AND2X1_RVT U594 ( .A1(n21), .A2(n65), .Y(ab_11__4_) );
  AND2X1_RVT U595 ( .A1(A[11]), .A2(n62), .Y(ab_11__3_) );
  AND2X1_RVT U596 ( .A1(n21), .A2(n61), .Y(ab_11__2_) );
  AND2X1_RVT U597 ( .A1(A[11]), .A2(n15), .Y(ab_11__20_) );
  AND2X1_RVT U598 ( .A1(n21), .A2(n59), .Y(ab_11__1_) );
  AND2X1_RVT U599 ( .A1(A[11]), .A2(n14), .Y(ab_11__19_) );
  AND2X1_RVT U600 ( .A1(n21), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U601 ( .A1(n21), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U602 ( .A1(n21), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U603 ( .A1(n21), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U604 ( .A1(n21), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U605 ( .A1(n21), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U606 ( .A1(n21), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U607 ( .A1(n21), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U608 ( .A1(n21), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U609 ( .A1(A[11]), .A2(n57), .Y(ab_11__0_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n75), .Y(ab_10__9_) );
  AND2X1_RVT U611 ( .A1(n20), .A2(n73), .Y(ab_10__8_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n71), .Y(ab_10__7_) );
  AND2X1_RVT U613 ( .A1(n20), .A2(n69), .Y(ab_10__6_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n67), .Y(ab_10__5_) );
  AND2X1_RVT U615 ( .A1(n20), .A2(n65), .Y(ab_10__4_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n63), .Y(ab_10__3_) );
  AND2X1_RVT U617 ( .A1(n20), .A2(n61), .Y(ab_10__2_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n16), .Y(ab_10__21_) );
  AND2X1_RVT U619 ( .A1(n20), .A2(n15), .Y(ab_10__20_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n59), .Y(ab_10__1_) );
  AND2X1_RVT U621 ( .A1(n20), .A2(n14), .Y(ab_10__19_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U623 ( .A1(n20), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U625 ( .A1(n20), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U627 ( .A1(n20), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U629 ( .A1(n20), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U631 ( .A1(n20), .A2(n57), .Y(ab_10__0_) );
  AND2X1_RVT U632 ( .A1(n36), .A2(n75), .Y(ab_0__9_) );
  AND2X1_RVT U633 ( .A1(n36), .A2(n73), .Y(ab_0__8_) );
  AND2X1_RVT U634 ( .A1(n36), .A2(n71), .Y(ab_0__7_) );
  AND2X1_RVT U635 ( .A1(n36), .A2(n69), .Y(ab_0__6_) );
  AND2X1_RVT U636 ( .A1(n36), .A2(n67), .Y(ab_0__5_) );
  AND2X1_RVT U637 ( .A1(n36), .A2(n64), .Y(ab_0__4_) );
  AND2X1_RVT U638 ( .A1(n36), .A2(n63), .Y(ab_0__3_) );
  AND2X1_RVT U639 ( .A1(n36), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U640 ( .A1(n35), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U641 ( .A1(n35), .A2(n61), .Y(ab_0__2_) );
  AND2X1_RVT U642 ( .A1(n35), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U643 ( .A1(n35), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U644 ( .A1(n35), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U645 ( .A1(n35), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U646 ( .A1(n35), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U647 ( .A1(n35), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U648 ( .A1(n35), .A2(n18), .Y(ab_0__23_) );
  AND2X1_RVT U649 ( .A1(n35), .A2(n17), .Y(ab_0__22_) );
  AND2X1_RVT U650 ( .A1(n35), .A2(n16), .Y(ab_0__21_) );
  AND2X1_RVT U651 ( .A1(n35), .A2(n15), .Y(ab_0__20_) );
  AND2X1_RVT U652 ( .A1(n34), .A2(n59), .Y(ab_0__1_) );
  AND2X1_RVT U653 ( .A1(n34), .A2(n14), .Y(ab_0__19_) );
  AND2X1_RVT U654 ( .A1(n34), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U655 ( .A1(n34), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U656 ( .A1(n34), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U657 ( .A1(n34), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U658 ( .A1(n34), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U659 ( .A1(n34), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U660 ( .A1(n34), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U661 ( .A1(n34), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U662 ( .A1(n34), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U663 ( .A1(n34), .A2(n57), .Y(PRODUCT_0_) );
endmodule


module OSPE_13_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_13 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n2), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n3), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n4), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n4), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n4), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n4), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n4), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n4), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n2), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n3), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n4), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n1), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n1), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n1), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n1), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n1), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n1), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n1), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n1), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n1), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n1), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n1), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n1), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n1), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n1), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n2), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n2), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n2), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n2), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n2), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n2), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n2), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n2), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n2), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n2), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n2), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n2), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_13_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_13_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_12_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n54) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n57) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n56) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n53) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n59) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n61) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n55) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n58) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n60) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n40) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n52) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n50) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n74) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n48) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n73) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n41) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n33) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n46) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n63) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n65) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n67) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n70) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n69) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n51) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n47) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n49) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n43) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n45) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n72) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n71) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n42) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n39) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n37) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n35) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n44) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n62) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n34) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n64) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n36) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n66) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n38) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n68) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n51), .A2(n74), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n49), .A2(n74), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n47), .A2(n74), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n45), .A2(n74), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n43), .A2(n74), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n41), .A2(n74), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n40), .A2(n74), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n38), .A2(n74), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n74), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n74), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n74), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n36), .A2(n73), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n73), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n73), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n73), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n73), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n73), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n73), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n73), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n73), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n73), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n73), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n33), .A2(n73), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n72), .A2(n51), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n72), .A2(n49), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n72), .A2(n47), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n72), .A2(n45), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n72), .A2(n43), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n72), .A2(n41), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n72), .A2(n40), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n72), .A2(n38), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n72), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n72), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n72), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n72), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n71), .A2(n36), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n71), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n71), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n71), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n71), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n71), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n71), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n71), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n71), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n71), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n71), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n71), .A2(n33), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n69), .A2(n51), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n70), .A2(n49), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n70), .A2(n47), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n70), .A2(n45), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n70), .A2(n43), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n70), .A2(n41), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n70), .A2(n40), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n70), .A2(n38), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n70), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n70), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n70), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n70), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n70), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n69), .A2(n36), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n69), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n69), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n69), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n69), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n69), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n69), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n69), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n69), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n69), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n69), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n69), .A2(n33), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n68), .A2(n51), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n68), .A2(n49), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n67), .A2(n47), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n67), .A2(n45), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n67), .A2(n43), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n67), .A2(n41), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n67), .A2(n40), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n67), .A2(n38), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n67), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n67), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n67), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n67), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n67), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n67), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n68), .A2(n36), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n68), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n68), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n68), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n68), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n68), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n68), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n68), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n68), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n68), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n68), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n68), .A2(n33), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n66), .A2(n51), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n66), .A2(n49), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n66), .A2(n47), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n65), .A2(n45), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n65), .A2(n43), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n65), .A2(n41), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n65), .A2(n40), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n65), .A2(n38), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n65), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n65), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n65), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n65), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n65), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n65), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n65), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n66), .A2(n36), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n66), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n66), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n66), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n66), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n66), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n66), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n66), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n66), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n66), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n66), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n66), .A2(n33), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n64), .A2(n51), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n64), .A2(n49), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n64), .A2(n47), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n64), .A2(n45), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n63), .A2(n43), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n63), .A2(n41), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n63), .A2(n40), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n63), .A2(n38), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n63), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n63), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n63), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n63), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n63), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n63), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n63), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n63), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n64), .A2(n36), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n64), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n64), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n64), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n64), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n64), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n64), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n64), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n64), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n64), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n64), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n64), .A2(n33), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n62), .A2(n51), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n62), .A2(n49), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n62), .A2(n47), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n62), .A2(n45), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n62), .A2(n43), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n61), .A2(n41), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n61), .A2(n40), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n61), .A2(n38), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n61), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n61), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n61), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n61), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n61), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n61), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n61), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n61), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n61), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n62), .A2(n36), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n62), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n62), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n62), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n62), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n62), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n62), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n62), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n62), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n62), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n62), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n62), .A2(n33), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n33), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n36), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n33), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n60), .A2(n51), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n60), .A2(n49), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n60), .A2(n47), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n60), .A2(n45), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n60), .A2(n43), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n60), .A2(n41), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n60), .A2(n40), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n59), .A2(n38), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n60), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n59), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n59), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n59), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n60), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n59), .A2(n36), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n59), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n59), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n59), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n59), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n59), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n59), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n59), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n59), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n59), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n59), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n59), .A2(n33), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n38), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n36), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n33), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n40), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n38), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n36), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n33), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n41), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n40), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n38), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n36), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n33), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n43), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n41), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n40), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n38), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n36), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n34), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n45), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n43), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n41), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n40), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n38), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n35), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n34), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n47), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n45), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n43), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n41), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n40), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n37), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n35), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n34), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n49), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n47), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n45), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n43), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n41), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n39), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n37), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n35), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n34), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n51), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n49), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n47), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n45), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n43), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n42), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n39), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n37), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n35), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n34), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n51), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n49), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n47), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n45), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n44), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n42), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n39), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n37), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n35), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n34), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n51), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n49), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n47), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n46), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n44), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n42), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n39), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n37), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n35), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n34), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n58), .A2(n51), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n58), .A2(n49), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n58), .A2(n48), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n58), .A2(n46), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n58), .A2(n44), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n58), .A2(n42), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n58), .A2(n39), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n57), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n57), .A2(n37), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n57), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n57), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n57), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n57), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n57), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n57), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n57), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n57), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n57), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n57), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n56), .A2(n35), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n56), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n56), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n56), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n56), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n56), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n56), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n56), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n56), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n56), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n56), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n56), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n51), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n50), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n48), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n46), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n44), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n42), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n39), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n37), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n35), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n34), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n52), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n50), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n48), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n46), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n44), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n42), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n39), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n37), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n35), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n34), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n52), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n50), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n48), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n46), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n44), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n42), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n39), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n37), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n35), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n34), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n52), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n50), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n48), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n46), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n44), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n42), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n39), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n37), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n35), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n34), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n52), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n50), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n48), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n46), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n44), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n42), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n39), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n37), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n35), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n34), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n52), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n50), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n48), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n46), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n44), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n42), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n39), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n37), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n35), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n34), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n52), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n50), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n48), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n46), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n44), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n42), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n39), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n37), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n35), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n34), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n52), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n50), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n48), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n46), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n44), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n42), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n39), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n37), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n36), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n34), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n52), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n50), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n48), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n46), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n44), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n42), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n39), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n38), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n36), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n34), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n52), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n50), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n48), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n46), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n44), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n42), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n40), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n38), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n36), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n34), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n55), .A2(n52), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n55), .A2(n50), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n55), .A2(n48), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n55), .A2(n46), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n55), .A2(n44), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n55), .A2(n41), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n55), .A2(n40), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n55), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n54), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n54), .A2(n38), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n54), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n54), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n54), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n54), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n54), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n54), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n54), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n54), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n54), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n54), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n53), .A2(n36), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n53), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n53), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n53), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n53), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n53), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n53), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n53), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n53), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n53), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n53), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n53), .A2(n34), .Y(PRODUCT_0_) );
endmodule


module OSPE_12_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_12 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n2), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n4), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n4), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n3), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n4), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n4), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n4), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n4), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n4), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n3), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n2), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n1), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n1), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n1), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n1), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n1), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n1), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n1), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n1), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n1), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n1), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n1), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n1), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n1), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n1), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n2), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n2), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n2), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n2), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n2), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n2), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n2), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n2), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n2), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n2), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n2), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n2), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_12_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_12_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_11_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_11_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_11 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n2), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n4), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n4), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n3), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n4), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n4), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n4), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n4), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n4), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n3), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n2), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n1), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n1), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n1), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n1), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n1), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n1), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n1), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n1), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n1), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n1), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n1), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n1), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n1), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n1), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n2), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n2), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n2), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n2), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n2), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n2), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n2), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n2), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n2), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n2), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n2), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n2), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_11_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_11_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_10_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U7 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U8 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U9 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U10 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U11 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U12 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U13 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U14 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_10_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_10 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n3), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n2), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n1), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n3), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n2), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n1), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n1), .Y(N100) );
  OSPE_10_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_10_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_9_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_9_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_9 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n1), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n2), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n1), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n2), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n1), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_9_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_9_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_8_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U4 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U5 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U6 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U7 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U8 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U9 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U10 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U11 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U12 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U13 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U14 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR2X1_RVT U15 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U16 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U17 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U18 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U19 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U20 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U21 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U22 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n53) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n56) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n55) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n52) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n58) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n60) );
  NBUFFX2_RVT U29 ( .A(A[4]), .Y(n62) );
  XOR2X1_RVT U30 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U31 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U32 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U33 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U34 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U35 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U36 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U37 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U38 ( .A(A[0]), .Y(n54) );
  NBUFFX2_RVT U39 ( .A(A[1]), .Y(n57) );
  XOR2X1_RVT U40 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U41 ( .A(A[2]), .Y(n59) );
  NBUFFX2_RVT U42 ( .A(B[3]), .Y(n39) );
  NBUFFX2_RVT U43 ( .A(A[9]), .Y(n73) );
  NBUFFX2_RVT U44 ( .A(B[9]), .Y(n51) );
  NBUFFX2_RVT U45 ( .A(A[9]), .Y(n72) );
  NBUFFX2_RVT U46 ( .A(B[8]), .Y(n49) );
  NBUFFX2_RVT U47 ( .A(A[5]), .Y(n64) );
  NBUFFX2_RVT U48 ( .A(A[6]), .Y(n66) );
  NBUFFX2_RVT U49 ( .A(A[7]), .Y(n69) );
  NBUFFX2_RVT U50 ( .A(A[7]), .Y(n68) );
  NBUFFX2_RVT U51 ( .A(B[7]), .Y(n47) );
  NBUFFX2_RVT U52 ( .A(A[8]), .Y(n71) );
  NBUFFX2_RVT U53 ( .A(A[8]), .Y(n70) );
  NBUFFX2_RVT U54 ( .A(B[4]), .Y(n40) );
  NBUFFX2_RVT U55 ( .A(B[0]), .Y(n32) );
  NBUFFX2_RVT U56 ( .A(B[6]), .Y(n45) );
  NBUFFX2_RVT U57 ( .A(B[9]), .Y(n50) );
  NBUFFX2_RVT U58 ( .A(B[7]), .Y(n46) );
  NBUFFX2_RVT U59 ( .A(B[8]), .Y(n48) );
  NBUFFX2_RVT U60 ( .A(B[5]), .Y(n42) );
  NBUFFX2_RVT U61 ( .A(B[6]), .Y(n44) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n41) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n38) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n36) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n34) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n43) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n61) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n33) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n63) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n35) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n65) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n37) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n67) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  NBUFFX2_RVT U131 ( .A(A[20]), .Y(n29) );
  NBUFFX2_RVT U132 ( .A(A[21]), .Y(n30) );
  NBUFFX2_RVT U133 ( .A(A[22]), .Y(n31) );
  AND2X1_RVT U134 ( .A1(n50), .A2(n73), .Y(ab_9__9_) );
  AND2X1_RVT U135 ( .A1(n48), .A2(n73), .Y(ab_9__8_) );
  AND2X1_RVT U136 ( .A1(n46), .A2(n73), .Y(ab_9__7_) );
  AND2X1_RVT U137 ( .A1(n44), .A2(n73), .Y(ab_9__6_) );
  AND2X1_RVT U138 ( .A1(n42), .A2(n73), .Y(ab_9__5_) );
  AND2X1_RVT U139 ( .A1(n40), .A2(n73), .Y(ab_9__4_) );
  AND2X1_RVT U140 ( .A1(n39), .A2(n73), .Y(ab_9__3_) );
  AND2X1_RVT U141 ( .A1(n37), .A2(n73), .Y(ab_9__2_) );
  AND2X1_RVT U142 ( .A1(B[22]), .A2(n73), .Y(ab_9__22_) );
  AND2X1_RVT U143 ( .A1(B[21]), .A2(n73), .Y(ab_9__21_) );
  AND2X1_RVT U144 ( .A1(n17), .A2(n73), .Y(ab_9__20_) );
  AND2X1_RVT U145 ( .A1(n35), .A2(n72), .Y(ab_9__1_) );
  AND2X1_RVT U146 ( .A1(n15), .A2(n72), .Y(ab_9__19_) );
  AND2X1_RVT U147 ( .A1(n13), .A2(n72), .Y(ab_9__18_) );
  AND2X1_RVT U148 ( .A1(B[17]), .A2(n72), .Y(ab_9__17_) );
  AND2X1_RVT U149 ( .A1(n11), .A2(n72), .Y(ab_9__16_) );
  AND2X1_RVT U150 ( .A1(n10), .A2(n72), .Y(ab_9__15_) );
  AND2X1_RVT U151 ( .A1(n9), .A2(n72), .Y(ab_9__14_) );
  AND2X1_RVT U152 ( .A1(B[13]), .A2(n72), .Y(ab_9__13_) );
  AND2X1_RVT U153 ( .A1(n7), .A2(n72), .Y(ab_9__12_) );
  AND2X1_RVT U154 ( .A1(n5), .A2(n72), .Y(ab_9__11_) );
  AND2X1_RVT U155 ( .A1(n3), .A2(n72), .Y(ab_9__10_) );
  AND2X1_RVT U156 ( .A1(n32), .A2(n72), .Y(ab_9__0_) );
  AND2X1_RVT U157 ( .A1(n71), .A2(n50), .Y(ab_8__9_) );
  AND2X1_RVT U158 ( .A1(n71), .A2(n48), .Y(ab_8__8_) );
  AND2X1_RVT U159 ( .A1(n71), .A2(n46), .Y(ab_8__7_) );
  AND2X1_RVT U160 ( .A1(n71), .A2(n44), .Y(ab_8__6_) );
  AND2X1_RVT U161 ( .A1(n71), .A2(n42), .Y(ab_8__5_) );
  AND2X1_RVT U162 ( .A1(n71), .A2(n40), .Y(ab_8__4_) );
  AND2X1_RVT U163 ( .A1(n71), .A2(n39), .Y(ab_8__3_) );
  AND2X1_RVT U164 ( .A1(n71), .A2(n37), .Y(ab_8__2_) );
  AND2X1_RVT U165 ( .A1(n71), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U166 ( .A1(n71), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U167 ( .A1(n71), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U168 ( .A1(n71), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U169 ( .A1(n70), .A2(n35), .Y(ab_8__1_) );
  AND2X1_RVT U170 ( .A1(n70), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U171 ( .A1(n70), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U172 ( .A1(n70), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U173 ( .A1(n70), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U174 ( .A1(n70), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U175 ( .A1(n70), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U176 ( .A1(n70), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U177 ( .A1(n70), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U178 ( .A1(n70), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U179 ( .A1(n70), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U180 ( .A1(n70), .A2(n32), .Y(ab_8__0_) );
  AND2X1_RVT U181 ( .A1(n68), .A2(n50), .Y(ab_7__9_) );
  AND2X1_RVT U182 ( .A1(n69), .A2(n48), .Y(ab_7__8_) );
  AND2X1_RVT U183 ( .A1(n69), .A2(n46), .Y(ab_7__7_) );
  AND2X1_RVT U184 ( .A1(n69), .A2(n44), .Y(ab_7__6_) );
  AND2X1_RVT U185 ( .A1(n69), .A2(n42), .Y(ab_7__5_) );
  AND2X1_RVT U186 ( .A1(n69), .A2(n40), .Y(ab_7__4_) );
  AND2X1_RVT U187 ( .A1(n69), .A2(n39), .Y(ab_7__3_) );
  AND2X1_RVT U188 ( .A1(n69), .A2(n37), .Y(ab_7__2_) );
  AND2X1_RVT U189 ( .A1(n69), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U190 ( .A1(n69), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U191 ( .A1(n69), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U192 ( .A1(n69), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U193 ( .A1(n69), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U194 ( .A1(n68), .A2(n35), .Y(ab_7__1_) );
  AND2X1_RVT U195 ( .A1(n68), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U196 ( .A1(n68), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U197 ( .A1(n68), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U198 ( .A1(n68), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U199 ( .A1(n68), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U200 ( .A1(n68), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U201 ( .A1(n68), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U202 ( .A1(n68), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U203 ( .A1(n68), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U204 ( .A1(n68), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U205 ( .A1(n68), .A2(n32), .Y(ab_7__0_) );
  AND2X1_RVT U206 ( .A1(n67), .A2(n50), .Y(ab_6__9_) );
  AND2X1_RVT U207 ( .A1(n67), .A2(n48), .Y(ab_6__8_) );
  AND2X1_RVT U208 ( .A1(n66), .A2(n46), .Y(ab_6__7_) );
  AND2X1_RVT U209 ( .A1(n66), .A2(n44), .Y(ab_6__6_) );
  AND2X1_RVT U210 ( .A1(n66), .A2(n42), .Y(ab_6__5_) );
  AND2X1_RVT U211 ( .A1(n66), .A2(n40), .Y(ab_6__4_) );
  AND2X1_RVT U212 ( .A1(n66), .A2(n39), .Y(ab_6__3_) );
  AND2X1_RVT U213 ( .A1(n66), .A2(n37), .Y(ab_6__2_) );
  AND2X1_RVT U214 ( .A1(n66), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U215 ( .A1(n66), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U216 ( .A1(n66), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U217 ( .A1(n66), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U218 ( .A1(n66), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U219 ( .A1(n66), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U220 ( .A1(n67), .A2(n35), .Y(ab_6__1_) );
  AND2X1_RVT U221 ( .A1(n67), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U222 ( .A1(n67), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U223 ( .A1(n67), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U224 ( .A1(n67), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U225 ( .A1(n67), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U226 ( .A1(n67), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U227 ( .A1(n67), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U228 ( .A1(n67), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U229 ( .A1(n67), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U230 ( .A1(n67), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U231 ( .A1(n67), .A2(n32), .Y(ab_6__0_) );
  AND2X1_RVT U232 ( .A1(n65), .A2(n50), .Y(ab_5__9_) );
  AND2X1_RVT U233 ( .A1(n65), .A2(n48), .Y(ab_5__8_) );
  AND2X1_RVT U234 ( .A1(n65), .A2(n46), .Y(ab_5__7_) );
  AND2X1_RVT U235 ( .A1(n64), .A2(n44), .Y(ab_5__6_) );
  AND2X1_RVT U236 ( .A1(n64), .A2(n42), .Y(ab_5__5_) );
  AND2X1_RVT U237 ( .A1(n64), .A2(n40), .Y(ab_5__4_) );
  AND2X1_RVT U238 ( .A1(n64), .A2(n39), .Y(ab_5__3_) );
  AND2X1_RVT U239 ( .A1(n64), .A2(n37), .Y(ab_5__2_) );
  AND2X1_RVT U240 ( .A1(n64), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U241 ( .A1(n64), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U242 ( .A1(n64), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U243 ( .A1(n64), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U244 ( .A1(n64), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U245 ( .A1(n64), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U246 ( .A1(n64), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U247 ( .A1(n65), .A2(n35), .Y(ab_5__1_) );
  AND2X1_RVT U248 ( .A1(n65), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U249 ( .A1(n65), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U250 ( .A1(n65), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U251 ( .A1(n65), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U252 ( .A1(n65), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U253 ( .A1(n65), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U254 ( .A1(n65), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U255 ( .A1(n65), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U256 ( .A1(n65), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U257 ( .A1(n65), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U258 ( .A1(n65), .A2(n32), .Y(ab_5__0_) );
  AND2X1_RVT U259 ( .A1(n63), .A2(n50), .Y(ab_4__9_) );
  AND2X1_RVT U260 ( .A1(n63), .A2(n48), .Y(ab_4__8_) );
  AND2X1_RVT U261 ( .A1(n63), .A2(n46), .Y(ab_4__7_) );
  AND2X1_RVT U262 ( .A1(n63), .A2(n44), .Y(ab_4__6_) );
  AND2X1_RVT U263 ( .A1(n62), .A2(n42), .Y(ab_4__5_) );
  AND2X1_RVT U264 ( .A1(n62), .A2(n40), .Y(ab_4__4_) );
  AND2X1_RVT U265 ( .A1(n62), .A2(n39), .Y(ab_4__3_) );
  AND2X1_RVT U266 ( .A1(n62), .A2(n37), .Y(ab_4__2_) );
  AND2X1_RVT U267 ( .A1(n62), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U268 ( .A1(n62), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U269 ( .A1(n62), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U270 ( .A1(n62), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U271 ( .A1(n62), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U272 ( .A1(n62), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U273 ( .A1(n62), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U274 ( .A1(n62), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U275 ( .A1(n63), .A2(n35), .Y(ab_4__1_) );
  AND2X1_RVT U276 ( .A1(n63), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U277 ( .A1(n63), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U278 ( .A1(n63), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U279 ( .A1(n63), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U280 ( .A1(n63), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U281 ( .A1(n63), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U282 ( .A1(n63), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U283 ( .A1(n63), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U284 ( .A1(n63), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U285 ( .A1(n63), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U286 ( .A1(n63), .A2(n32), .Y(ab_4__0_) );
  AND2X1_RVT U287 ( .A1(n61), .A2(n50), .Y(ab_3__9_) );
  AND2X1_RVT U288 ( .A1(n61), .A2(n48), .Y(ab_3__8_) );
  AND2X1_RVT U289 ( .A1(n61), .A2(n46), .Y(ab_3__7_) );
  AND2X1_RVT U290 ( .A1(n61), .A2(n44), .Y(ab_3__6_) );
  AND2X1_RVT U291 ( .A1(n61), .A2(n42), .Y(ab_3__5_) );
  AND2X1_RVT U292 ( .A1(n60), .A2(n40), .Y(ab_3__4_) );
  AND2X1_RVT U293 ( .A1(n60), .A2(n39), .Y(ab_3__3_) );
  AND2X1_RVT U294 ( .A1(n60), .A2(n37), .Y(ab_3__2_) );
  AND2X1_RVT U295 ( .A1(n60), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U296 ( .A1(n60), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U297 ( .A1(n60), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U298 ( .A1(n60), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U299 ( .A1(n60), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U300 ( .A1(n60), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U301 ( .A1(n60), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U302 ( .A1(n60), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U303 ( .A1(n60), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U304 ( .A1(n61), .A2(n35), .Y(ab_3__1_) );
  AND2X1_RVT U305 ( .A1(n61), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U306 ( .A1(n61), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U307 ( .A1(n61), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U308 ( .A1(n61), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U309 ( .A1(n61), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U310 ( .A1(n61), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U311 ( .A1(n61), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U312 ( .A1(n61), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U313 ( .A1(n61), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U314 ( .A1(n61), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U315 ( .A1(n61), .A2(n32), .Y(ab_3__0_) );
  AND2X1_RVT U316 ( .A1(A[31]), .A2(n32), .Y(ab_31__0_) );
  AND2X1_RVT U317 ( .A1(A[30]), .A2(n35), .Y(ab_30__1_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n32), .Y(ab_30__0_) );
  AND2X1_RVT U319 ( .A1(n59), .A2(n50), .Y(ab_2__9_) );
  AND2X1_RVT U320 ( .A1(n59), .A2(n48), .Y(ab_2__8_) );
  AND2X1_RVT U321 ( .A1(n59), .A2(n46), .Y(ab_2__7_) );
  AND2X1_RVT U322 ( .A1(n59), .A2(n44), .Y(ab_2__6_) );
  AND2X1_RVT U323 ( .A1(n59), .A2(n42), .Y(ab_2__5_) );
  AND2X1_RVT U324 ( .A1(n59), .A2(n40), .Y(ab_2__4_) );
  AND2X1_RVT U325 ( .A1(n59), .A2(n39), .Y(ab_2__3_) );
  AND2X1_RVT U326 ( .A1(n58), .A2(n37), .Y(ab_2__2_) );
  AND2X1_RVT U327 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U329 ( .A1(n59), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U330 ( .A1(n58), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U331 ( .A1(n58), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U332 ( .A1(n58), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U333 ( .A1(n59), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U335 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U337 ( .A1(n58), .A2(n35), .Y(ab_2__1_) );
  AND2X1_RVT U338 ( .A1(n58), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U339 ( .A1(n58), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U340 ( .A1(n58), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U341 ( .A1(n58), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U342 ( .A1(n58), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U343 ( .A1(n58), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U344 ( .A1(n58), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U345 ( .A1(n58), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U346 ( .A1(n58), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U347 ( .A1(n58), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U348 ( .A1(n58), .A2(n32), .Y(ab_2__0_) );
  AND2X1_RVT U349 ( .A1(A[29]), .A2(n37), .Y(ab_29__2_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n35), .Y(ab_29__1_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n32), .Y(ab_29__0_) );
  AND2X1_RVT U352 ( .A1(A[28]), .A2(n39), .Y(ab_28__3_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n37), .Y(ab_28__2_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n35), .Y(ab_28__1_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n32), .Y(ab_28__0_) );
  AND2X1_RVT U356 ( .A1(A[27]), .A2(n40), .Y(ab_27__4_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n39), .Y(ab_27__3_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n37), .Y(ab_27__2_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n35), .Y(ab_27__1_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n32), .Y(ab_27__0_) );
  AND2X1_RVT U361 ( .A1(A[26]), .A2(n42), .Y(ab_26__5_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n40), .Y(ab_26__4_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n39), .Y(ab_26__3_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n37), .Y(ab_26__2_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n35), .Y(ab_26__1_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n33), .Y(ab_26__0_) );
  AND2X1_RVT U367 ( .A1(A[25]), .A2(n44), .Y(ab_25__6_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n42), .Y(ab_25__5_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n40), .Y(ab_25__4_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n39), .Y(ab_25__3_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n37), .Y(ab_25__2_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n34), .Y(ab_25__1_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n33), .Y(ab_25__0_) );
  AND2X1_RVT U374 ( .A1(A[24]), .A2(n46), .Y(ab_24__7_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n44), .Y(ab_24__6_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n42), .Y(ab_24__5_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n40), .Y(ab_24__4_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n39), .Y(ab_24__3_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n36), .Y(ab_24__2_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n34), .Y(ab_24__1_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n33), .Y(ab_24__0_) );
  AND2X1_RVT U382 ( .A1(A[23]), .A2(n48), .Y(ab_23__8_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n46), .Y(ab_23__7_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n44), .Y(ab_23__6_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n42), .Y(ab_23__5_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n40), .Y(ab_23__4_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n38), .Y(ab_23__3_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n36), .Y(ab_23__2_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n34), .Y(ab_23__1_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n33), .Y(ab_23__0_) );
  AND2X1_RVT U391 ( .A1(A[22]), .A2(n50), .Y(ab_22__9_) );
  AND2X1_RVT U392 ( .A1(n31), .A2(n48), .Y(ab_22__8_) );
  AND2X1_RVT U393 ( .A1(n31), .A2(n46), .Y(ab_22__7_) );
  AND2X1_RVT U394 ( .A1(n31), .A2(n44), .Y(ab_22__6_) );
  AND2X1_RVT U395 ( .A1(n31), .A2(n42), .Y(ab_22__5_) );
  AND2X1_RVT U396 ( .A1(n31), .A2(n41), .Y(ab_22__4_) );
  AND2X1_RVT U397 ( .A1(n31), .A2(n38), .Y(ab_22__3_) );
  AND2X1_RVT U398 ( .A1(n31), .A2(n36), .Y(ab_22__2_) );
  AND2X1_RVT U399 ( .A1(n31), .A2(n34), .Y(ab_22__1_) );
  AND2X1_RVT U400 ( .A1(n31), .A2(n33), .Y(ab_22__0_) );
  AND2X1_RVT U401 ( .A1(n30), .A2(n50), .Y(ab_21__9_) );
  AND2X1_RVT U402 ( .A1(n30), .A2(n48), .Y(ab_21__8_) );
  AND2X1_RVT U403 ( .A1(n30), .A2(n46), .Y(ab_21__7_) );
  AND2X1_RVT U404 ( .A1(n30), .A2(n44), .Y(ab_21__6_) );
  AND2X1_RVT U405 ( .A1(n30), .A2(n43), .Y(ab_21__5_) );
  AND2X1_RVT U406 ( .A1(n30), .A2(n41), .Y(ab_21__4_) );
  AND2X1_RVT U407 ( .A1(n30), .A2(n38), .Y(ab_21__3_) );
  AND2X1_RVT U408 ( .A1(n30), .A2(n36), .Y(ab_21__2_) );
  AND2X1_RVT U409 ( .A1(n30), .A2(n34), .Y(ab_21__1_) );
  AND2X1_RVT U410 ( .A1(n30), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U411 ( .A1(n30), .A2(n33), .Y(ab_21__0_) );
  AND2X1_RVT U412 ( .A1(n29), .A2(n50), .Y(ab_20__9_) );
  AND2X1_RVT U413 ( .A1(n29), .A2(n48), .Y(ab_20__8_) );
  AND2X1_RVT U414 ( .A1(n29), .A2(n46), .Y(ab_20__7_) );
  AND2X1_RVT U415 ( .A1(n29), .A2(n45), .Y(ab_20__6_) );
  AND2X1_RVT U416 ( .A1(n29), .A2(n43), .Y(ab_20__5_) );
  AND2X1_RVT U417 ( .A1(n29), .A2(n41), .Y(ab_20__4_) );
  AND2X1_RVT U418 ( .A1(n29), .A2(n38), .Y(ab_20__3_) );
  AND2X1_RVT U419 ( .A1(n29), .A2(n36), .Y(ab_20__2_) );
  AND2X1_RVT U420 ( .A1(n29), .A2(n34), .Y(ab_20__1_) );
  AND2X1_RVT U421 ( .A1(n29), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U422 ( .A1(n29), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U423 ( .A1(n29), .A2(n33), .Y(ab_20__0_) );
  AND2X1_RVT U424 ( .A1(n57), .A2(n50), .Y(ab_1__9_) );
  AND2X1_RVT U425 ( .A1(n57), .A2(n48), .Y(ab_1__8_) );
  AND2X1_RVT U426 ( .A1(n57), .A2(n47), .Y(ab_1__7_) );
  AND2X1_RVT U427 ( .A1(n57), .A2(n45), .Y(ab_1__6_) );
  AND2X1_RVT U428 ( .A1(n57), .A2(n43), .Y(ab_1__5_) );
  AND2X1_RVT U429 ( .A1(n57), .A2(n41), .Y(ab_1__4_) );
  AND2X1_RVT U430 ( .A1(n57), .A2(n38), .Y(ab_1__3_) );
  AND2X1_RVT U431 ( .A1(n56), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U432 ( .A1(n56), .A2(n36), .Y(ab_1__2_) );
  AND2X1_RVT U433 ( .A1(n56), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U434 ( .A1(n56), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U435 ( .A1(n56), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U436 ( .A1(n56), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U437 ( .A1(n56), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U438 ( .A1(n56), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U439 ( .A1(n56), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U440 ( .A1(n56), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U441 ( .A1(n56), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U442 ( .A1(n56), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U443 ( .A1(n55), .A2(n34), .Y(ab_1__1_) );
  AND2X1_RVT U444 ( .A1(n55), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U445 ( .A1(n55), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U446 ( .A1(n55), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U447 ( .A1(n55), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U448 ( .A1(n55), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U449 ( .A1(n55), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U450 ( .A1(n55), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U451 ( .A1(n55), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U452 ( .A1(n55), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U453 ( .A1(n55), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U454 ( .A1(n55), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U455 ( .A1(n28), .A2(n50), .Y(ab_19__9_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n49), .Y(ab_19__8_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n47), .Y(ab_19__7_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n45), .Y(ab_19__6_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n43), .Y(ab_19__5_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n41), .Y(ab_19__4_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n38), .Y(ab_19__3_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n36), .Y(ab_19__2_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n34), .Y(ab_19__1_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U467 ( .A1(A[19]), .A2(n33), .Y(ab_19__0_) );
  AND2X1_RVT U468 ( .A1(n27), .A2(n51), .Y(ab_18__9_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n49), .Y(ab_18__8_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n47), .Y(ab_18__7_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n45), .Y(ab_18__6_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n43), .Y(ab_18__5_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n41), .Y(ab_18__4_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n38), .Y(ab_18__3_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n36), .Y(ab_18__2_) );
  AND2X1_RVT U476 ( .A1(A[18]), .A2(n34), .Y(ab_18__1_) );
  AND2X1_RVT U477 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n33), .Y(ab_18__0_) );
  AND2X1_RVT U482 ( .A1(n26), .A2(n51), .Y(ab_17__9_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n49), .Y(ab_17__8_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n47), .Y(ab_17__7_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n45), .Y(ab_17__6_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n43), .Y(ab_17__5_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n41), .Y(ab_17__4_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n38), .Y(ab_17__3_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n36), .Y(ab_17__2_) );
  AND2X1_RVT U490 ( .A1(A[17]), .A2(n34), .Y(ab_17__1_) );
  AND2X1_RVT U491 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U496 ( .A1(A[17]), .A2(n33), .Y(ab_17__0_) );
  AND2X1_RVT U497 ( .A1(n25), .A2(n51), .Y(ab_16__9_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n49), .Y(ab_16__8_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n47), .Y(ab_16__7_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n45), .Y(ab_16__6_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n43), .Y(ab_16__5_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n41), .Y(ab_16__4_) );
  AND2X1_RVT U503 ( .A1(A[16]), .A2(n38), .Y(ab_16__3_) );
  AND2X1_RVT U504 ( .A1(n25), .A2(n36), .Y(ab_16__2_) );
  AND2X1_RVT U505 ( .A1(A[16]), .A2(n34), .Y(ab_16__1_) );
  AND2X1_RVT U506 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n33), .Y(ab_16__0_) );
  AND2X1_RVT U513 ( .A1(n24), .A2(n51), .Y(ab_15__9_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n49), .Y(ab_15__8_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n47), .Y(ab_15__7_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n45), .Y(ab_15__6_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n43), .Y(ab_15__5_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n41), .Y(ab_15__4_) );
  AND2X1_RVT U519 ( .A1(A[15]), .A2(n38), .Y(ab_15__3_) );
  AND2X1_RVT U520 ( .A1(n24), .A2(n36), .Y(ab_15__2_) );
  AND2X1_RVT U521 ( .A1(A[15]), .A2(n34), .Y(ab_15__1_) );
  AND2X1_RVT U522 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U529 ( .A1(A[15]), .A2(n33), .Y(ab_15__0_) );
  AND2X1_RVT U530 ( .A1(n23), .A2(n51), .Y(ab_14__9_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n49), .Y(ab_14__8_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n47), .Y(ab_14__7_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n45), .Y(ab_14__6_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n43), .Y(ab_14__5_) );
  AND2X1_RVT U535 ( .A1(A[14]), .A2(n41), .Y(ab_14__4_) );
  AND2X1_RVT U536 ( .A1(n23), .A2(n38), .Y(ab_14__3_) );
  AND2X1_RVT U537 ( .A1(A[14]), .A2(n36), .Y(ab_14__2_) );
  AND2X1_RVT U538 ( .A1(n23), .A2(n34), .Y(ab_14__1_) );
  AND2X1_RVT U539 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U540 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U547 ( .A1(A[14]), .A2(n33), .Y(ab_14__0_) );
  AND2X1_RVT U548 ( .A1(n22), .A2(n51), .Y(ab_13__9_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n49), .Y(ab_13__8_) );
  AND2X1_RVT U550 ( .A1(A[13]), .A2(n47), .Y(ab_13__7_) );
  AND2X1_RVT U551 ( .A1(n22), .A2(n45), .Y(ab_13__6_) );
  AND2X1_RVT U552 ( .A1(A[13]), .A2(n43), .Y(ab_13__5_) );
  AND2X1_RVT U553 ( .A1(n22), .A2(n41), .Y(ab_13__4_) );
  AND2X1_RVT U554 ( .A1(A[13]), .A2(n38), .Y(ab_13__3_) );
  AND2X1_RVT U555 ( .A1(n22), .A2(n36), .Y(ab_13__2_) );
  AND2X1_RVT U556 ( .A1(A[13]), .A2(n34), .Y(ab_13__1_) );
  AND2X1_RVT U557 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U566 ( .A1(A[13]), .A2(n33), .Y(ab_13__0_) );
  AND2X1_RVT U567 ( .A1(n21), .A2(n51), .Y(ab_12__9_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n49), .Y(ab_12__8_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n47), .Y(ab_12__7_) );
  AND2X1_RVT U570 ( .A1(A[12]), .A2(n45), .Y(ab_12__6_) );
  AND2X1_RVT U571 ( .A1(n21), .A2(n43), .Y(ab_12__5_) );
  AND2X1_RVT U572 ( .A1(A[12]), .A2(n41), .Y(ab_12__4_) );
  AND2X1_RVT U573 ( .A1(n21), .A2(n38), .Y(ab_12__3_) );
  AND2X1_RVT U574 ( .A1(A[12]), .A2(n36), .Y(ab_12__2_) );
  AND2X1_RVT U575 ( .A1(n21), .A2(n35), .Y(ab_12__1_) );
  AND2X1_RVT U576 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U577 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U586 ( .A1(A[12]), .A2(n33), .Y(ab_12__0_) );
  AND2X1_RVT U587 ( .A1(n20), .A2(n51), .Y(ab_11__9_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n49), .Y(ab_11__8_) );
  AND2X1_RVT U589 ( .A1(A[11]), .A2(n47), .Y(ab_11__7_) );
  AND2X1_RVT U590 ( .A1(n20), .A2(n45), .Y(ab_11__6_) );
  AND2X1_RVT U591 ( .A1(A[11]), .A2(n43), .Y(ab_11__5_) );
  AND2X1_RVT U592 ( .A1(n20), .A2(n41), .Y(ab_11__4_) );
  AND2X1_RVT U593 ( .A1(A[11]), .A2(n38), .Y(ab_11__3_) );
  AND2X1_RVT U594 ( .A1(n20), .A2(n37), .Y(ab_11__2_) );
  AND2X1_RVT U595 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U596 ( .A1(n20), .A2(n35), .Y(ab_11__1_) );
  AND2X1_RVT U597 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U598 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U607 ( .A1(A[11]), .A2(n33), .Y(ab_11__0_) );
  AND2X1_RVT U608 ( .A1(n18), .A2(n51), .Y(ab_10__9_) );
  AND2X1_RVT U609 ( .A1(n19), .A2(n49), .Y(ab_10__8_) );
  AND2X1_RVT U610 ( .A1(n18), .A2(n47), .Y(ab_10__7_) );
  AND2X1_RVT U611 ( .A1(n19), .A2(n45), .Y(ab_10__6_) );
  AND2X1_RVT U612 ( .A1(n18), .A2(n43), .Y(ab_10__5_) );
  AND2X1_RVT U613 ( .A1(n19), .A2(n41), .Y(ab_10__4_) );
  AND2X1_RVT U614 ( .A1(n18), .A2(n39), .Y(ab_10__3_) );
  AND2X1_RVT U615 ( .A1(n19), .A2(n37), .Y(ab_10__2_) );
  AND2X1_RVT U616 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U617 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U618 ( .A1(n18), .A2(n35), .Y(ab_10__1_) );
  AND2X1_RVT U619 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U620 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U621 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U622 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U623 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U624 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U625 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U626 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U627 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U628 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U629 ( .A1(n19), .A2(n33), .Y(ab_10__0_) );
  AND2X1_RVT U630 ( .A1(n54), .A2(n51), .Y(ab_0__9_) );
  AND2X1_RVT U631 ( .A1(n54), .A2(n49), .Y(ab_0__8_) );
  AND2X1_RVT U632 ( .A1(n54), .A2(n47), .Y(ab_0__7_) );
  AND2X1_RVT U633 ( .A1(n54), .A2(n45), .Y(ab_0__6_) );
  AND2X1_RVT U634 ( .A1(n54), .A2(n43), .Y(ab_0__5_) );
  AND2X1_RVT U635 ( .A1(n54), .A2(n40), .Y(ab_0__4_) );
  AND2X1_RVT U636 ( .A1(n54), .A2(n39), .Y(ab_0__3_) );
  AND2X1_RVT U637 ( .A1(n54), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U638 ( .A1(n53), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U639 ( .A1(n53), .A2(n37), .Y(ab_0__2_) );
  AND2X1_RVT U640 ( .A1(n53), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U641 ( .A1(n53), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U642 ( .A1(n53), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U643 ( .A1(n53), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U644 ( .A1(n53), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U645 ( .A1(n53), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U646 ( .A1(n53), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U647 ( .A1(n53), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U648 ( .A1(n53), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U649 ( .A1(n53), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U650 ( .A1(n52), .A2(n35), .Y(ab_0__1_) );
  AND2X1_RVT U651 ( .A1(n52), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U652 ( .A1(n52), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U653 ( .A1(n52), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U654 ( .A1(n52), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U655 ( .A1(n52), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U656 ( .A1(n52), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U657 ( .A1(n52), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U658 ( .A1(n52), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U659 ( .A1(n52), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U660 ( .A1(n52), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U661 ( .A1(n52), .A2(n33), .Y(PRODUCT_0_) );
endmodule


module OSPE_8_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_8 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n1), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n3), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n2), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n1), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n3), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n2), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n1), .Y(N100) );
  OSPE_8_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_8_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_7_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_7_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_7 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n1), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n2), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n1), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n2), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n1), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_7_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_7_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_6_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U7 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U8 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U9 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U10 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U11 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U12 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U13 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U14 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U15 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U16 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U17 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_6_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_6 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n1), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n3), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n2), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n1), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n3), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n2), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n1), .Y(N100) );
  OSPE_6_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_6_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_5_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_5_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_5 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n3), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n2), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n4), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n3), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n2), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n4), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n4), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n4), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n4), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n4), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n4), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n1), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n1), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n1), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n1), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n1), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n1), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n1), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n1), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n1), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n1), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n1), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n1), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n1), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n1), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n2), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n2), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n2), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n2), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n2), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n2), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n2), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n2), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n2), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n2), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n2), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n2), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n2), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n2), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n3), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n3), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n3), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n3), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n3), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n3), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n3), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n3), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n3), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n3), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n3), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n3), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n3), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n3), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n4), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n4), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n4), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n4), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n4), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n4), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n5), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n5), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n6), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n6), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n6), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n6), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n6), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n6), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n6), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n6), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n5), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n5), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n5), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n5), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n5), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n5), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n5), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n5), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n5), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n5), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n5), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n5), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n5), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n5), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n6), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n6), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n6), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n6), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n6), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n4), .Y(N100) );
  OSPE_5_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_5_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
endmodule


module OSPE_4_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U4 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U5 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U6 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U7 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U8 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U9 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U10 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U11 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U12 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U13 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U14 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  XOR2X1_RVT U15 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U16 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U17 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U18 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U19 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U20 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U21 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U22 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n53) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n56) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n55) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n52) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n58) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n60) );
  NBUFFX2_RVT U29 ( .A(A[4]), .Y(n62) );
  XOR2X1_RVT U30 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U31 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U32 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U33 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U34 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U35 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U36 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U37 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U38 ( .A(A[0]), .Y(n54) );
  NBUFFX2_RVT U39 ( .A(A[1]), .Y(n57) );
  XOR2X1_RVT U40 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U41 ( .A(A[2]), .Y(n59) );
  NBUFFX2_RVT U42 ( .A(B[3]), .Y(n39) );
  NBUFFX2_RVT U43 ( .A(A[9]), .Y(n73) );
  NBUFFX2_RVT U44 ( .A(B[9]), .Y(n51) );
  NBUFFX2_RVT U45 ( .A(A[9]), .Y(n72) );
  NBUFFX2_RVT U46 ( .A(B[8]), .Y(n49) );
  NBUFFX2_RVT U47 ( .A(A[5]), .Y(n64) );
  NBUFFX2_RVT U48 ( .A(A[6]), .Y(n66) );
  NBUFFX2_RVT U49 ( .A(A[7]), .Y(n69) );
  NBUFFX2_RVT U50 ( .A(A[7]), .Y(n68) );
  NBUFFX2_RVT U51 ( .A(B[7]), .Y(n47) );
  NBUFFX2_RVT U52 ( .A(A[8]), .Y(n71) );
  NBUFFX2_RVT U53 ( .A(A[8]), .Y(n70) );
  NBUFFX2_RVT U54 ( .A(B[4]), .Y(n40) );
  NBUFFX2_RVT U55 ( .A(B[0]), .Y(n32) );
  NBUFFX2_RVT U56 ( .A(B[6]), .Y(n45) );
  NBUFFX2_RVT U57 ( .A(B[9]), .Y(n50) );
  NBUFFX2_RVT U58 ( .A(B[7]), .Y(n46) );
  NBUFFX2_RVT U59 ( .A(B[8]), .Y(n48) );
  NBUFFX2_RVT U60 ( .A(B[5]), .Y(n42) );
  NBUFFX2_RVT U61 ( .A(B[6]), .Y(n44) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n41) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n38) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n36) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n34) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n43) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n61) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n33) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n63) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n35) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n65) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n37) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n67) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  NBUFFX2_RVT U131 ( .A(A[20]), .Y(n29) );
  NBUFFX2_RVT U132 ( .A(A[21]), .Y(n30) );
  NBUFFX2_RVT U133 ( .A(A[22]), .Y(n31) );
  AND2X1_RVT U134 ( .A1(n50), .A2(n73), .Y(ab_9__9_) );
  AND2X1_RVT U135 ( .A1(n48), .A2(n73), .Y(ab_9__8_) );
  AND2X1_RVT U136 ( .A1(n46), .A2(n73), .Y(ab_9__7_) );
  AND2X1_RVT U137 ( .A1(n44), .A2(n73), .Y(ab_9__6_) );
  AND2X1_RVT U138 ( .A1(n42), .A2(n73), .Y(ab_9__5_) );
  AND2X1_RVT U139 ( .A1(n40), .A2(n73), .Y(ab_9__4_) );
  AND2X1_RVT U140 ( .A1(n39), .A2(n73), .Y(ab_9__3_) );
  AND2X1_RVT U141 ( .A1(n37), .A2(n73), .Y(ab_9__2_) );
  AND2X1_RVT U142 ( .A1(B[22]), .A2(n73), .Y(ab_9__22_) );
  AND2X1_RVT U143 ( .A1(B[21]), .A2(n73), .Y(ab_9__21_) );
  AND2X1_RVT U144 ( .A1(n17), .A2(n73), .Y(ab_9__20_) );
  AND2X1_RVT U145 ( .A1(n35), .A2(n72), .Y(ab_9__1_) );
  AND2X1_RVT U146 ( .A1(n15), .A2(n72), .Y(ab_9__19_) );
  AND2X1_RVT U147 ( .A1(n13), .A2(n72), .Y(ab_9__18_) );
  AND2X1_RVT U148 ( .A1(B[17]), .A2(n72), .Y(ab_9__17_) );
  AND2X1_RVT U149 ( .A1(n11), .A2(n72), .Y(ab_9__16_) );
  AND2X1_RVT U150 ( .A1(n10), .A2(n72), .Y(ab_9__15_) );
  AND2X1_RVT U151 ( .A1(n9), .A2(n72), .Y(ab_9__14_) );
  AND2X1_RVT U152 ( .A1(B[13]), .A2(n72), .Y(ab_9__13_) );
  AND2X1_RVT U153 ( .A1(n7), .A2(n72), .Y(ab_9__12_) );
  AND2X1_RVT U154 ( .A1(n5), .A2(n72), .Y(ab_9__11_) );
  AND2X1_RVT U155 ( .A1(n3), .A2(n72), .Y(ab_9__10_) );
  AND2X1_RVT U156 ( .A1(n32), .A2(n72), .Y(ab_9__0_) );
  AND2X1_RVT U157 ( .A1(n71), .A2(n50), .Y(ab_8__9_) );
  AND2X1_RVT U158 ( .A1(n71), .A2(n48), .Y(ab_8__8_) );
  AND2X1_RVT U159 ( .A1(n71), .A2(n46), .Y(ab_8__7_) );
  AND2X1_RVT U160 ( .A1(n71), .A2(n44), .Y(ab_8__6_) );
  AND2X1_RVT U161 ( .A1(n71), .A2(n42), .Y(ab_8__5_) );
  AND2X1_RVT U162 ( .A1(n71), .A2(n40), .Y(ab_8__4_) );
  AND2X1_RVT U163 ( .A1(n71), .A2(n39), .Y(ab_8__3_) );
  AND2X1_RVT U164 ( .A1(n71), .A2(n37), .Y(ab_8__2_) );
  AND2X1_RVT U165 ( .A1(n71), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U166 ( .A1(n71), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U167 ( .A1(n71), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U168 ( .A1(n71), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U169 ( .A1(n70), .A2(n35), .Y(ab_8__1_) );
  AND2X1_RVT U170 ( .A1(n70), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U171 ( .A1(n70), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U172 ( .A1(n70), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U173 ( .A1(n70), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U174 ( .A1(n70), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U175 ( .A1(n70), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U176 ( .A1(n70), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U177 ( .A1(n70), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U178 ( .A1(n70), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U179 ( .A1(n70), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U180 ( .A1(n70), .A2(n32), .Y(ab_8__0_) );
  AND2X1_RVT U181 ( .A1(n68), .A2(n50), .Y(ab_7__9_) );
  AND2X1_RVT U182 ( .A1(n69), .A2(n48), .Y(ab_7__8_) );
  AND2X1_RVT U183 ( .A1(n69), .A2(n46), .Y(ab_7__7_) );
  AND2X1_RVT U184 ( .A1(n69), .A2(n44), .Y(ab_7__6_) );
  AND2X1_RVT U185 ( .A1(n69), .A2(n42), .Y(ab_7__5_) );
  AND2X1_RVT U186 ( .A1(n69), .A2(n40), .Y(ab_7__4_) );
  AND2X1_RVT U187 ( .A1(n69), .A2(n39), .Y(ab_7__3_) );
  AND2X1_RVT U188 ( .A1(n69), .A2(n37), .Y(ab_7__2_) );
  AND2X1_RVT U189 ( .A1(n69), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U190 ( .A1(n69), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U191 ( .A1(n69), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U192 ( .A1(n69), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U193 ( .A1(n69), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U194 ( .A1(n68), .A2(n35), .Y(ab_7__1_) );
  AND2X1_RVT U195 ( .A1(n68), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U196 ( .A1(n68), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U197 ( .A1(n68), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U198 ( .A1(n68), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U199 ( .A1(n68), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U200 ( .A1(n68), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U201 ( .A1(n68), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U202 ( .A1(n68), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U203 ( .A1(n68), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U204 ( .A1(n68), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U205 ( .A1(n68), .A2(n32), .Y(ab_7__0_) );
  AND2X1_RVT U206 ( .A1(n67), .A2(n50), .Y(ab_6__9_) );
  AND2X1_RVT U207 ( .A1(n67), .A2(n48), .Y(ab_6__8_) );
  AND2X1_RVT U208 ( .A1(n66), .A2(n46), .Y(ab_6__7_) );
  AND2X1_RVT U209 ( .A1(n66), .A2(n44), .Y(ab_6__6_) );
  AND2X1_RVT U210 ( .A1(n66), .A2(n42), .Y(ab_6__5_) );
  AND2X1_RVT U211 ( .A1(n66), .A2(n40), .Y(ab_6__4_) );
  AND2X1_RVT U212 ( .A1(n66), .A2(n39), .Y(ab_6__3_) );
  AND2X1_RVT U213 ( .A1(n66), .A2(n37), .Y(ab_6__2_) );
  AND2X1_RVT U214 ( .A1(n66), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U215 ( .A1(n66), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U216 ( .A1(n66), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U217 ( .A1(n66), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U218 ( .A1(n66), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U219 ( .A1(n66), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U220 ( .A1(n67), .A2(n35), .Y(ab_6__1_) );
  AND2X1_RVT U221 ( .A1(n67), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U222 ( .A1(n67), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U223 ( .A1(n67), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U224 ( .A1(n67), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U225 ( .A1(n67), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U226 ( .A1(n67), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U227 ( .A1(n67), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U228 ( .A1(n67), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U229 ( .A1(n67), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U230 ( .A1(n67), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U231 ( .A1(n67), .A2(n32), .Y(ab_6__0_) );
  AND2X1_RVT U232 ( .A1(n65), .A2(n50), .Y(ab_5__9_) );
  AND2X1_RVT U233 ( .A1(n65), .A2(n48), .Y(ab_5__8_) );
  AND2X1_RVT U234 ( .A1(n65), .A2(n46), .Y(ab_5__7_) );
  AND2X1_RVT U235 ( .A1(n64), .A2(n44), .Y(ab_5__6_) );
  AND2X1_RVT U236 ( .A1(n64), .A2(n42), .Y(ab_5__5_) );
  AND2X1_RVT U237 ( .A1(n64), .A2(n40), .Y(ab_5__4_) );
  AND2X1_RVT U238 ( .A1(n64), .A2(n39), .Y(ab_5__3_) );
  AND2X1_RVT U239 ( .A1(n64), .A2(n37), .Y(ab_5__2_) );
  AND2X1_RVT U240 ( .A1(n64), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U241 ( .A1(n64), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U242 ( .A1(n64), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U243 ( .A1(n64), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U244 ( .A1(n64), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U245 ( .A1(n64), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U246 ( .A1(n64), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U247 ( .A1(n65), .A2(n35), .Y(ab_5__1_) );
  AND2X1_RVT U248 ( .A1(n65), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U249 ( .A1(n65), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U250 ( .A1(n65), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U251 ( .A1(n65), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U252 ( .A1(n65), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U253 ( .A1(n65), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U254 ( .A1(n65), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U255 ( .A1(n65), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U256 ( .A1(n65), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U257 ( .A1(n65), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U258 ( .A1(n65), .A2(n32), .Y(ab_5__0_) );
  AND2X1_RVT U259 ( .A1(n63), .A2(n50), .Y(ab_4__9_) );
  AND2X1_RVT U260 ( .A1(n63), .A2(n48), .Y(ab_4__8_) );
  AND2X1_RVT U261 ( .A1(n63), .A2(n46), .Y(ab_4__7_) );
  AND2X1_RVT U262 ( .A1(n63), .A2(n44), .Y(ab_4__6_) );
  AND2X1_RVT U263 ( .A1(n62), .A2(n42), .Y(ab_4__5_) );
  AND2X1_RVT U264 ( .A1(n62), .A2(n40), .Y(ab_4__4_) );
  AND2X1_RVT U265 ( .A1(n62), .A2(n39), .Y(ab_4__3_) );
  AND2X1_RVT U266 ( .A1(n62), .A2(n37), .Y(ab_4__2_) );
  AND2X1_RVT U267 ( .A1(n62), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U268 ( .A1(n62), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U269 ( .A1(n62), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U270 ( .A1(n62), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U271 ( .A1(n62), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U272 ( .A1(n62), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U273 ( .A1(n62), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U274 ( .A1(n62), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U275 ( .A1(n63), .A2(n35), .Y(ab_4__1_) );
  AND2X1_RVT U276 ( .A1(n63), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U277 ( .A1(n63), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U278 ( .A1(n63), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U279 ( .A1(n63), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U280 ( .A1(n63), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U281 ( .A1(n63), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U282 ( .A1(n63), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U283 ( .A1(n63), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U284 ( .A1(n63), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U285 ( .A1(n63), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U286 ( .A1(n63), .A2(n32), .Y(ab_4__0_) );
  AND2X1_RVT U287 ( .A1(n61), .A2(n50), .Y(ab_3__9_) );
  AND2X1_RVT U288 ( .A1(n61), .A2(n48), .Y(ab_3__8_) );
  AND2X1_RVT U289 ( .A1(n61), .A2(n46), .Y(ab_3__7_) );
  AND2X1_RVT U290 ( .A1(n61), .A2(n44), .Y(ab_3__6_) );
  AND2X1_RVT U291 ( .A1(n61), .A2(n42), .Y(ab_3__5_) );
  AND2X1_RVT U292 ( .A1(n60), .A2(n40), .Y(ab_3__4_) );
  AND2X1_RVT U293 ( .A1(n60), .A2(n39), .Y(ab_3__3_) );
  AND2X1_RVT U294 ( .A1(n60), .A2(n37), .Y(ab_3__2_) );
  AND2X1_RVT U295 ( .A1(n60), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U296 ( .A1(n60), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U297 ( .A1(n60), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U298 ( .A1(n60), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U299 ( .A1(n60), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U300 ( .A1(n60), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U301 ( .A1(n60), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U302 ( .A1(n60), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U303 ( .A1(n60), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U304 ( .A1(n61), .A2(n35), .Y(ab_3__1_) );
  AND2X1_RVT U305 ( .A1(n61), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U306 ( .A1(n61), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U307 ( .A1(n61), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U308 ( .A1(n61), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U309 ( .A1(n61), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U310 ( .A1(n61), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U311 ( .A1(n61), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U312 ( .A1(n61), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U313 ( .A1(n61), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U314 ( .A1(n61), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U315 ( .A1(n61), .A2(n32), .Y(ab_3__0_) );
  AND2X1_RVT U316 ( .A1(A[31]), .A2(n32), .Y(ab_31__0_) );
  AND2X1_RVT U317 ( .A1(A[30]), .A2(n35), .Y(ab_30__1_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n32), .Y(ab_30__0_) );
  AND2X1_RVT U319 ( .A1(n59), .A2(n50), .Y(ab_2__9_) );
  AND2X1_RVT U320 ( .A1(n59), .A2(n48), .Y(ab_2__8_) );
  AND2X1_RVT U321 ( .A1(n59), .A2(n46), .Y(ab_2__7_) );
  AND2X1_RVT U322 ( .A1(n59), .A2(n44), .Y(ab_2__6_) );
  AND2X1_RVT U323 ( .A1(n59), .A2(n42), .Y(ab_2__5_) );
  AND2X1_RVT U324 ( .A1(n59), .A2(n40), .Y(ab_2__4_) );
  AND2X1_RVT U325 ( .A1(n59), .A2(n39), .Y(ab_2__3_) );
  AND2X1_RVT U326 ( .A1(n58), .A2(n37), .Y(ab_2__2_) );
  AND2X1_RVT U327 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U329 ( .A1(n59), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U330 ( .A1(n58), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U331 ( .A1(n58), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U332 ( .A1(n58), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U333 ( .A1(n59), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U335 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U337 ( .A1(n58), .A2(n35), .Y(ab_2__1_) );
  AND2X1_RVT U338 ( .A1(n58), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U339 ( .A1(n58), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U340 ( .A1(n58), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U341 ( .A1(n58), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U342 ( .A1(n58), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U343 ( .A1(n58), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U344 ( .A1(n58), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U345 ( .A1(n58), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U346 ( .A1(n58), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U347 ( .A1(n58), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U348 ( .A1(n58), .A2(n32), .Y(ab_2__0_) );
  AND2X1_RVT U349 ( .A1(A[29]), .A2(n37), .Y(ab_29__2_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n35), .Y(ab_29__1_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n32), .Y(ab_29__0_) );
  AND2X1_RVT U352 ( .A1(A[28]), .A2(n39), .Y(ab_28__3_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n37), .Y(ab_28__2_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n35), .Y(ab_28__1_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n32), .Y(ab_28__0_) );
  AND2X1_RVT U356 ( .A1(A[27]), .A2(n40), .Y(ab_27__4_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n39), .Y(ab_27__3_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n37), .Y(ab_27__2_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n35), .Y(ab_27__1_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n32), .Y(ab_27__0_) );
  AND2X1_RVT U361 ( .A1(A[26]), .A2(n42), .Y(ab_26__5_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n40), .Y(ab_26__4_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n39), .Y(ab_26__3_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n37), .Y(ab_26__2_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n35), .Y(ab_26__1_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n33), .Y(ab_26__0_) );
  AND2X1_RVT U367 ( .A1(A[25]), .A2(n44), .Y(ab_25__6_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n42), .Y(ab_25__5_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n40), .Y(ab_25__4_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n39), .Y(ab_25__3_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n37), .Y(ab_25__2_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n34), .Y(ab_25__1_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n33), .Y(ab_25__0_) );
  AND2X1_RVT U374 ( .A1(A[24]), .A2(n46), .Y(ab_24__7_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n44), .Y(ab_24__6_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n42), .Y(ab_24__5_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n40), .Y(ab_24__4_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n39), .Y(ab_24__3_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n36), .Y(ab_24__2_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n34), .Y(ab_24__1_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n33), .Y(ab_24__0_) );
  AND2X1_RVT U382 ( .A1(A[23]), .A2(n48), .Y(ab_23__8_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n46), .Y(ab_23__7_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n44), .Y(ab_23__6_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n42), .Y(ab_23__5_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n40), .Y(ab_23__4_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n38), .Y(ab_23__3_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n36), .Y(ab_23__2_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n34), .Y(ab_23__1_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n33), .Y(ab_23__0_) );
  AND2X1_RVT U391 ( .A1(A[22]), .A2(n50), .Y(ab_22__9_) );
  AND2X1_RVT U392 ( .A1(n31), .A2(n48), .Y(ab_22__8_) );
  AND2X1_RVT U393 ( .A1(n31), .A2(n46), .Y(ab_22__7_) );
  AND2X1_RVT U394 ( .A1(n31), .A2(n44), .Y(ab_22__6_) );
  AND2X1_RVT U395 ( .A1(n31), .A2(n42), .Y(ab_22__5_) );
  AND2X1_RVT U396 ( .A1(n31), .A2(n41), .Y(ab_22__4_) );
  AND2X1_RVT U397 ( .A1(n31), .A2(n38), .Y(ab_22__3_) );
  AND2X1_RVT U398 ( .A1(n31), .A2(n36), .Y(ab_22__2_) );
  AND2X1_RVT U399 ( .A1(n31), .A2(n34), .Y(ab_22__1_) );
  AND2X1_RVT U400 ( .A1(n31), .A2(n33), .Y(ab_22__0_) );
  AND2X1_RVT U401 ( .A1(n30), .A2(n50), .Y(ab_21__9_) );
  AND2X1_RVT U402 ( .A1(n30), .A2(n48), .Y(ab_21__8_) );
  AND2X1_RVT U403 ( .A1(n30), .A2(n46), .Y(ab_21__7_) );
  AND2X1_RVT U404 ( .A1(n30), .A2(n44), .Y(ab_21__6_) );
  AND2X1_RVT U405 ( .A1(n30), .A2(n43), .Y(ab_21__5_) );
  AND2X1_RVT U406 ( .A1(n30), .A2(n41), .Y(ab_21__4_) );
  AND2X1_RVT U407 ( .A1(n30), .A2(n38), .Y(ab_21__3_) );
  AND2X1_RVT U408 ( .A1(n30), .A2(n36), .Y(ab_21__2_) );
  AND2X1_RVT U409 ( .A1(n30), .A2(n34), .Y(ab_21__1_) );
  AND2X1_RVT U410 ( .A1(n30), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U411 ( .A1(n30), .A2(n33), .Y(ab_21__0_) );
  AND2X1_RVT U412 ( .A1(n29), .A2(n50), .Y(ab_20__9_) );
  AND2X1_RVT U413 ( .A1(n29), .A2(n48), .Y(ab_20__8_) );
  AND2X1_RVT U414 ( .A1(n29), .A2(n46), .Y(ab_20__7_) );
  AND2X1_RVT U415 ( .A1(n29), .A2(n45), .Y(ab_20__6_) );
  AND2X1_RVT U416 ( .A1(n29), .A2(n43), .Y(ab_20__5_) );
  AND2X1_RVT U417 ( .A1(n29), .A2(n41), .Y(ab_20__4_) );
  AND2X1_RVT U418 ( .A1(n29), .A2(n38), .Y(ab_20__3_) );
  AND2X1_RVT U419 ( .A1(n29), .A2(n36), .Y(ab_20__2_) );
  AND2X1_RVT U420 ( .A1(n29), .A2(n34), .Y(ab_20__1_) );
  AND2X1_RVT U421 ( .A1(n29), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U422 ( .A1(n29), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U423 ( .A1(n29), .A2(n33), .Y(ab_20__0_) );
  AND2X1_RVT U424 ( .A1(n57), .A2(n50), .Y(ab_1__9_) );
  AND2X1_RVT U425 ( .A1(n57), .A2(n48), .Y(ab_1__8_) );
  AND2X1_RVT U426 ( .A1(n57), .A2(n47), .Y(ab_1__7_) );
  AND2X1_RVT U427 ( .A1(n57), .A2(n45), .Y(ab_1__6_) );
  AND2X1_RVT U428 ( .A1(n57), .A2(n43), .Y(ab_1__5_) );
  AND2X1_RVT U429 ( .A1(n57), .A2(n41), .Y(ab_1__4_) );
  AND2X1_RVT U430 ( .A1(n57), .A2(n38), .Y(ab_1__3_) );
  AND2X1_RVT U431 ( .A1(n56), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U432 ( .A1(n56), .A2(n36), .Y(ab_1__2_) );
  AND2X1_RVT U433 ( .A1(n56), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U434 ( .A1(n56), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U435 ( .A1(n56), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U436 ( .A1(n56), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U437 ( .A1(n56), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U438 ( .A1(n56), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U439 ( .A1(n56), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U440 ( .A1(n56), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U441 ( .A1(n56), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U442 ( .A1(n56), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U443 ( .A1(n55), .A2(n34), .Y(ab_1__1_) );
  AND2X1_RVT U444 ( .A1(n55), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U445 ( .A1(n55), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U446 ( .A1(n55), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U447 ( .A1(n55), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U448 ( .A1(n55), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U449 ( .A1(n55), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U450 ( .A1(n55), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U451 ( .A1(n55), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U452 ( .A1(n55), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U453 ( .A1(n55), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U454 ( .A1(n55), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U455 ( .A1(n28), .A2(n50), .Y(ab_19__9_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n49), .Y(ab_19__8_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n47), .Y(ab_19__7_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n45), .Y(ab_19__6_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n43), .Y(ab_19__5_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n41), .Y(ab_19__4_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n38), .Y(ab_19__3_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n36), .Y(ab_19__2_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n34), .Y(ab_19__1_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U467 ( .A1(A[19]), .A2(n33), .Y(ab_19__0_) );
  AND2X1_RVT U468 ( .A1(n27), .A2(n51), .Y(ab_18__9_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n49), .Y(ab_18__8_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n47), .Y(ab_18__7_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n45), .Y(ab_18__6_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n43), .Y(ab_18__5_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n41), .Y(ab_18__4_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n38), .Y(ab_18__3_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n36), .Y(ab_18__2_) );
  AND2X1_RVT U476 ( .A1(A[18]), .A2(n34), .Y(ab_18__1_) );
  AND2X1_RVT U477 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n33), .Y(ab_18__0_) );
  AND2X1_RVT U482 ( .A1(n26), .A2(n51), .Y(ab_17__9_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n49), .Y(ab_17__8_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n47), .Y(ab_17__7_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n45), .Y(ab_17__6_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n43), .Y(ab_17__5_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n41), .Y(ab_17__4_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n38), .Y(ab_17__3_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n36), .Y(ab_17__2_) );
  AND2X1_RVT U490 ( .A1(A[17]), .A2(n34), .Y(ab_17__1_) );
  AND2X1_RVT U491 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U496 ( .A1(A[17]), .A2(n33), .Y(ab_17__0_) );
  AND2X1_RVT U497 ( .A1(n25), .A2(n51), .Y(ab_16__9_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n49), .Y(ab_16__8_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n47), .Y(ab_16__7_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n45), .Y(ab_16__6_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n43), .Y(ab_16__5_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n41), .Y(ab_16__4_) );
  AND2X1_RVT U503 ( .A1(A[16]), .A2(n38), .Y(ab_16__3_) );
  AND2X1_RVT U504 ( .A1(n25), .A2(n36), .Y(ab_16__2_) );
  AND2X1_RVT U505 ( .A1(A[16]), .A2(n34), .Y(ab_16__1_) );
  AND2X1_RVT U506 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n33), .Y(ab_16__0_) );
  AND2X1_RVT U513 ( .A1(n24), .A2(n51), .Y(ab_15__9_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n49), .Y(ab_15__8_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n47), .Y(ab_15__7_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n45), .Y(ab_15__6_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n43), .Y(ab_15__5_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n41), .Y(ab_15__4_) );
  AND2X1_RVT U519 ( .A1(A[15]), .A2(n38), .Y(ab_15__3_) );
  AND2X1_RVT U520 ( .A1(n24), .A2(n36), .Y(ab_15__2_) );
  AND2X1_RVT U521 ( .A1(A[15]), .A2(n34), .Y(ab_15__1_) );
  AND2X1_RVT U522 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U529 ( .A1(A[15]), .A2(n33), .Y(ab_15__0_) );
  AND2X1_RVT U530 ( .A1(n23), .A2(n51), .Y(ab_14__9_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n49), .Y(ab_14__8_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n47), .Y(ab_14__7_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n45), .Y(ab_14__6_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n43), .Y(ab_14__5_) );
  AND2X1_RVT U535 ( .A1(A[14]), .A2(n41), .Y(ab_14__4_) );
  AND2X1_RVT U536 ( .A1(n23), .A2(n38), .Y(ab_14__3_) );
  AND2X1_RVT U537 ( .A1(A[14]), .A2(n36), .Y(ab_14__2_) );
  AND2X1_RVT U538 ( .A1(n23), .A2(n34), .Y(ab_14__1_) );
  AND2X1_RVT U539 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U540 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U547 ( .A1(A[14]), .A2(n33), .Y(ab_14__0_) );
  AND2X1_RVT U548 ( .A1(n22), .A2(n51), .Y(ab_13__9_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n49), .Y(ab_13__8_) );
  AND2X1_RVT U550 ( .A1(A[13]), .A2(n47), .Y(ab_13__7_) );
  AND2X1_RVT U551 ( .A1(n22), .A2(n45), .Y(ab_13__6_) );
  AND2X1_RVT U552 ( .A1(A[13]), .A2(n43), .Y(ab_13__5_) );
  AND2X1_RVT U553 ( .A1(n22), .A2(n41), .Y(ab_13__4_) );
  AND2X1_RVT U554 ( .A1(A[13]), .A2(n38), .Y(ab_13__3_) );
  AND2X1_RVT U555 ( .A1(n22), .A2(n36), .Y(ab_13__2_) );
  AND2X1_RVT U556 ( .A1(A[13]), .A2(n34), .Y(ab_13__1_) );
  AND2X1_RVT U557 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U566 ( .A1(A[13]), .A2(n33), .Y(ab_13__0_) );
  AND2X1_RVT U567 ( .A1(n21), .A2(n51), .Y(ab_12__9_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n49), .Y(ab_12__8_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n47), .Y(ab_12__7_) );
  AND2X1_RVT U570 ( .A1(A[12]), .A2(n45), .Y(ab_12__6_) );
  AND2X1_RVT U571 ( .A1(n21), .A2(n43), .Y(ab_12__5_) );
  AND2X1_RVT U572 ( .A1(A[12]), .A2(n41), .Y(ab_12__4_) );
  AND2X1_RVT U573 ( .A1(n21), .A2(n38), .Y(ab_12__3_) );
  AND2X1_RVT U574 ( .A1(A[12]), .A2(n36), .Y(ab_12__2_) );
  AND2X1_RVT U575 ( .A1(n21), .A2(n35), .Y(ab_12__1_) );
  AND2X1_RVT U576 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U577 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U586 ( .A1(A[12]), .A2(n33), .Y(ab_12__0_) );
  AND2X1_RVT U587 ( .A1(n20), .A2(n51), .Y(ab_11__9_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n49), .Y(ab_11__8_) );
  AND2X1_RVT U589 ( .A1(A[11]), .A2(n47), .Y(ab_11__7_) );
  AND2X1_RVT U590 ( .A1(n20), .A2(n45), .Y(ab_11__6_) );
  AND2X1_RVT U591 ( .A1(A[11]), .A2(n43), .Y(ab_11__5_) );
  AND2X1_RVT U592 ( .A1(n20), .A2(n41), .Y(ab_11__4_) );
  AND2X1_RVT U593 ( .A1(A[11]), .A2(n38), .Y(ab_11__3_) );
  AND2X1_RVT U594 ( .A1(n20), .A2(n37), .Y(ab_11__2_) );
  AND2X1_RVT U595 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U596 ( .A1(n20), .A2(n35), .Y(ab_11__1_) );
  AND2X1_RVT U597 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U598 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U607 ( .A1(A[11]), .A2(n33), .Y(ab_11__0_) );
  AND2X1_RVT U608 ( .A1(n18), .A2(n51), .Y(ab_10__9_) );
  AND2X1_RVT U609 ( .A1(n19), .A2(n49), .Y(ab_10__8_) );
  AND2X1_RVT U610 ( .A1(n18), .A2(n47), .Y(ab_10__7_) );
  AND2X1_RVT U611 ( .A1(n19), .A2(n45), .Y(ab_10__6_) );
  AND2X1_RVT U612 ( .A1(n18), .A2(n43), .Y(ab_10__5_) );
  AND2X1_RVT U613 ( .A1(n19), .A2(n41), .Y(ab_10__4_) );
  AND2X1_RVT U614 ( .A1(n18), .A2(n39), .Y(ab_10__3_) );
  AND2X1_RVT U615 ( .A1(n19), .A2(n37), .Y(ab_10__2_) );
  AND2X1_RVT U616 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U617 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U618 ( .A1(n18), .A2(n35), .Y(ab_10__1_) );
  AND2X1_RVT U619 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U620 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U621 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U622 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U623 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U624 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U625 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U626 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U627 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U628 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U629 ( .A1(n19), .A2(n33), .Y(ab_10__0_) );
  AND2X1_RVT U630 ( .A1(n54), .A2(n51), .Y(ab_0__9_) );
  AND2X1_RVT U631 ( .A1(n54), .A2(n49), .Y(ab_0__8_) );
  AND2X1_RVT U632 ( .A1(n54), .A2(n47), .Y(ab_0__7_) );
  AND2X1_RVT U633 ( .A1(n54), .A2(n45), .Y(ab_0__6_) );
  AND2X1_RVT U634 ( .A1(n54), .A2(n43), .Y(ab_0__5_) );
  AND2X1_RVT U635 ( .A1(n54), .A2(n40), .Y(ab_0__4_) );
  AND2X1_RVT U636 ( .A1(n54), .A2(n39), .Y(ab_0__3_) );
  AND2X1_RVT U637 ( .A1(n54), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U638 ( .A1(n53), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U639 ( .A1(n53), .A2(n37), .Y(ab_0__2_) );
  AND2X1_RVT U640 ( .A1(n53), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U641 ( .A1(n53), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U642 ( .A1(n53), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U643 ( .A1(n53), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U644 ( .A1(n53), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U645 ( .A1(n53), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U646 ( .A1(n53), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U647 ( .A1(n53), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U648 ( .A1(n53), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U649 ( .A1(n53), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U650 ( .A1(n52), .A2(n35), .Y(ab_0__1_) );
  AND2X1_RVT U651 ( .A1(n52), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U652 ( .A1(n52), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U653 ( .A1(n52), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U654 ( .A1(n52), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U655 ( .A1(n52), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U656 ( .A1(n52), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U657 ( .A1(n52), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U658 ( .A1(n52), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U659 ( .A1(n52), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U660 ( .A1(n52), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U661 ( .A1(n52), .A2(n33), .Y(PRODUCT_0_) );
endmodule


module OSPE_4_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_4 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33, N32,
         N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18,
         N17, N16, N15, N14, N13, N12, N11, N10, n2, n3, n4, n5, n6, n7;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n2), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n2), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n2), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n2), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n2), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n2), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n2), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n2), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n2), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n2), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n2), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n2), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n2), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n3), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n3), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n3), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n3), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n3), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n3), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n3), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n3), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n3), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n3), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n3), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n3), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n3), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n3), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n4), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n4), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n4), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n4), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n4), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n4), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n4), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n4), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n4), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n4), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n4), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n4), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n4), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n4), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n5), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n5), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n5), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n5), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n5), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n5), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n5), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n5), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n5), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n5), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n5), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n5), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n5), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n2), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n4), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n3), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n5), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n2), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n4), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n3), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n5), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n7), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n6), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n7), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n6), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n7), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n6), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n7), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n7), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n7), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n7), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n7), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n7), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n7), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n6), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n6), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n6), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n6), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n6), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n6), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n6), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n6), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n6), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n6), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n6), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n6), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n6), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n6), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n7), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n7), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n7), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n7), .Y(N103) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n2), .Y(N100) );
  OSPE_4_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_4_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  DFFSSRX1_RVT opC_reg_0_ ( .D(opC_wire[0]), .SETB(1'b1), .RSTB(n7), .CLK(clk), 
        .Q(opC[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n5) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U103 ( .A(rstnPsum), .Y(n6) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n7) );
endmodule


module OSPE_3_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_3_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_3 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6,
         n7;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n5), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n5), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n5), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n5), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n5), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n5), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n5), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n5), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n6), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n7), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n6), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n7), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n7), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n7), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n7), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n7), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n7), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n7), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n7), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n7), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n7), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n6), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n6), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n6), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n6), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n6), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n6), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n6), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n6), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n6), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n6), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n6), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n6), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n6), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n6), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n7), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n7), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n7), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n7), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n7), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n5), .Y(N100) );
  OSPE_3_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_3_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPipe), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
  NBUFFX2_RVT U105 ( .A(rstnPsum), .Y(n7) );
endmodule


module OSPE_2_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(n39), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(n39), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(A[2]), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n40), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_2_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_2 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6,
         n7;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n5), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n5), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n5), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n5), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n5), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n5), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n5), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n5), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n6), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n7), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n6), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n7), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n7), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n7), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n7), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n7), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n7), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n7), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n7), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n7), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n7), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n6), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n6), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n6), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n6), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n6), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n6), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n6), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n6), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n6), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n6), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n6), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n6), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n6), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n6), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n7), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n7), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n7), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n7), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n7), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n5), .Y(N100) );
  OSPE_2_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_2_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPipe), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
  NBUFFX2_RVT U105 ( .A(rstnPsum), .Y(n7) );
endmodule


module OSPE_1_DW02_mult_0 ( A, B, PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, 
        PRODUCT_28_, PRODUCT_27_, PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, 
        PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, 
        PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, 
        PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, 
        PRODUCT_8_, PRODUCT_7_, PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, 
        PRODUCT_2_, PRODUCT_1_, PRODUCT_0_ );
  input [31:0] A;
  input [31:0] B;
  output PRODUCT_31_, PRODUCT_30_, PRODUCT_29_, PRODUCT_28_, PRODUCT_27_,
         PRODUCT_26_, PRODUCT_25_, PRODUCT_24_, PRODUCT_23_, PRODUCT_22_,
         PRODUCT_21_, PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_,
         PRODUCT_16_, PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_,
         PRODUCT_11_, PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_,
         PRODUCT_6_, PRODUCT_5_, PRODUCT_4_, PRODUCT_3_, PRODUCT_2_,
         PRODUCT_1_, PRODUCT_0_;
  wire   ab_31__0_, ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_,
         ab_27__2_, ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_,
         ab_26__2_, ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_,
         ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__8_, ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_,
         ab_23__2_, ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_,
         ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_,
         ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_,
         ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_, ab_15__11_,
         ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_, ab_15__5_,
         ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__13_, ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_,
         ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_, ab_12__11_,
         ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_, ab_12__5_,
         ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__20_,
         ab_11__19_, ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_,
         ab_11__14_, ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_,
         ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_,
         ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_, ab_10__20_, ab_10__19_,
         ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_,
         ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__26_, ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_,
         ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_,
         ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_,
         ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_,
         ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_,
         ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_, ab_1__27_,
         ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_, ab_1__21_,
         ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_,
         ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_,
         ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_, ab_0__28_,
         ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_,
         ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__29_,
         CARRYB_1__28_, CARRYB_1__27_, CARRYB_1__26_, CARRYB_1__25_,
         CARRYB_1__24_, CARRYB_1__23_, CARRYB_1__22_, CARRYB_1__21_,
         CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_, CARRYB_1__17_,
         CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_, CARRYB_1__13_,
         CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_, CARRYB_1__9_,
         CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_,
         SUMB_1__29_, SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_,
         SUMB_1__24_, SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_,
         SUMB_1__19_, SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_,
         SUMB_1__14_, SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_,
         SUMB_1__9_, SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_,
         CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_,
         CARRYB_28__0_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_,
         CARRYB_26__1_, CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_,
         CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_,
         CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_,
         CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_,
         CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_,
         CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_,
         SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_,
         SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_,
         SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_,
         SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_,
         SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_,
         SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_,
         SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;

  FADDX1_RVT S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .S(
        PRODUCT_31_) );
  FADDX1_RVT S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(PRODUCT_30_) );
  FADDX1_RVT S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .S(
        SUMB_30__1_) );
  FADDX1_RVT S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(PRODUCT_29_) );
  FADDX1_RVT S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  FADDX1_RVT S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .S(
        SUMB_29__2_) );
  FADDX1_RVT S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(PRODUCT_28_) );
  FADDX1_RVT S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  FADDX1_RVT S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  FADDX1_RVT S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .S(
        SUMB_28__3_) );
  FADDX1_RVT S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(PRODUCT_27_) );
  FADDX1_RVT S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  FADDX1_RVT S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  FADDX1_RVT S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  FADDX1_RVT S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .S(
        SUMB_27__4_) );
  FADDX1_RVT S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(PRODUCT_26_) );
  FADDX1_RVT S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  FADDX1_RVT S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  FADDX1_RVT S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  FADDX1_RVT S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  FADDX1_RVT S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .S(
        SUMB_26__5_) );
  FADDX1_RVT S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(PRODUCT_25_) );
  FADDX1_RVT S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  FADDX1_RVT S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  FADDX1_RVT S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  FADDX1_RVT S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  FADDX1_RVT S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  FADDX1_RVT S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .S(
        SUMB_25__6_) );
  FADDX1_RVT S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(PRODUCT_24_) );
  FADDX1_RVT S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  FADDX1_RVT S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  FADDX1_RVT S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  FADDX1_RVT S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  FADDX1_RVT S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  FADDX1_RVT S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  FADDX1_RVT S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .S(
        SUMB_24__7_) );
  FADDX1_RVT S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(PRODUCT_23_) );
  FADDX1_RVT S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  FADDX1_RVT S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  FADDX1_RVT S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  FADDX1_RVT S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  FADDX1_RVT S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  FADDX1_RVT S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  FADDX1_RVT S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  FADDX1_RVT S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .S(
        SUMB_23__8_) );
  FADDX1_RVT S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(PRODUCT_22_) );
  FADDX1_RVT S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  FADDX1_RVT S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  FADDX1_RVT S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  FADDX1_RVT S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  FADDX1_RVT S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  FADDX1_RVT S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  FADDX1_RVT S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  FADDX1_RVT S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  FADDX1_RVT S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .S(SUMB_22__9_) );
  FADDX1_RVT S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(PRODUCT_21_) );
  FADDX1_RVT S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  FADDX1_RVT S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  FADDX1_RVT S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  FADDX1_RVT S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  FADDX1_RVT S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  FADDX1_RVT S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  FADDX1_RVT S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  FADDX1_RVT S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  FADDX1_RVT S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  FADDX1_RVT S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), 
        .S(SUMB_21__10_) );
  FADDX1_RVT S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(PRODUCT_20_) );
  FADDX1_RVT S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  FADDX1_RVT S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  FADDX1_RVT S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  FADDX1_RVT S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  FADDX1_RVT S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  FADDX1_RVT S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  FADDX1_RVT S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  FADDX1_RVT S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  FADDX1_RVT S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  FADDX1_RVT S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  FADDX1_RVT S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), 
        .S(SUMB_20__11_) );
  FADDX1_RVT S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(PRODUCT_19_) );
  FADDX1_RVT S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  FADDX1_RVT S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  FADDX1_RVT S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  FADDX1_RVT S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  FADDX1_RVT S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  FADDX1_RVT S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  FADDX1_RVT S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  FADDX1_RVT S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  FADDX1_RVT S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  FADDX1_RVT S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  FADDX1_RVT S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  FADDX1_RVT S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), 
        .S(SUMB_19__12_) );
  FADDX1_RVT S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(PRODUCT_18_) );
  FADDX1_RVT S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  FADDX1_RVT S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  FADDX1_RVT S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  FADDX1_RVT S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  FADDX1_RVT S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  FADDX1_RVT S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  FADDX1_RVT S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  FADDX1_RVT S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  FADDX1_RVT S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  FADDX1_RVT S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  FADDX1_RVT S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  FADDX1_RVT S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  FADDX1_RVT S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), 
        .S(SUMB_18__13_) );
  FADDX1_RVT S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(PRODUCT_17_) );
  FADDX1_RVT S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  FADDX1_RVT S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  FADDX1_RVT S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  FADDX1_RVT S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  FADDX1_RVT S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  FADDX1_RVT S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  FADDX1_RVT S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  FADDX1_RVT S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  FADDX1_RVT S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  FADDX1_RVT S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  FADDX1_RVT S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  FADDX1_RVT S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  FADDX1_RVT S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  FADDX1_RVT S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), 
        .S(SUMB_17__14_) );
  FADDX1_RVT S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(PRODUCT_16_) );
  FADDX1_RVT S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  FADDX1_RVT S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  FADDX1_RVT S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  FADDX1_RVT S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  FADDX1_RVT S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  FADDX1_RVT S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  FADDX1_RVT S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  FADDX1_RVT S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  FADDX1_RVT S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  FADDX1_RVT S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  FADDX1_RVT S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  FADDX1_RVT S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  FADDX1_RVT S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  FADDX1_RVT S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  FADDX1_RVT S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), 
        .S(SUMB_16__15_) );
  FADDX1_RVT S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(PRODUCT_15_) );
  FADDX1_RVT S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  FADDX1_RVT S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  FADDX1_RVT S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  FADDX1_RVT S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  FADDX1_RVT S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  FADDX1_RVT S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  FADDX1_RVT S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  FADDX1_RVT S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  FADDX1_RVT S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  FADDX1_RVT S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  FADDX1_RVT S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  FADDX1_RVT S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  FADDX1_RVT S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  FADDX1_RVT S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  FADDX1_RVT S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), 
        .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  FADDX1_RVT S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), 
        .S(SUMB_15__16_) );
  FADDX1_RVT S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(PRODUCT_14_) );
  FADDX1_RVT S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  FADDX1_RVT S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  FADDX1_RVT S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  FADDX1_RVT S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  FADDX1_RVT S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  FADDX1_RVT S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  FADDX1_RVT S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  FADDX1_RVT S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  FADDX1_RVT S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  FADDX1_RVT S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  FADDX1_RVT S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  FADDX1_RVT S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  FADDX1_RVT S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  FADDX1_RVT S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), 
        .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  FADDX1_RVT S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  FADDX1_RVT S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  FADDX1_RVT S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), 
        .S(SUMB_14__17_) );
  FADDX1_RVT S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(PRODUCT_13_) );
  FADDX1_RVT S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  FADDX1_RVT S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  FADDX1_RVT S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  FADDX1_RVT S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  FADDX1_RVT S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  FADDX1_RVT S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  FADDX1_RVT S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  FADDX1_RVT S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  FADDX1_RVT S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  FADDX1_RVT S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  FADDX1_RVT S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  FADDX1_RVT S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  FADDX1_RVT S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), 
        .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  FADDX1_RVT S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  FADDX1_RVT S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  FADDX1_RVT S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  FADDX1_RVT S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  FADDX1_RVT S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), 
        .S(SUMB_13__18_) );
  FADDX1_RVT S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(PRODUCT_12_) );
  FADDX1_RVT S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  FADDX1_RVT S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  FADDX1_RVT S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  FADDX1_RVT S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  FADDX1_RVT S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  FADDX1_RVT S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  FADDX1_RVT S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  FADDX1_RVT S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  FADDX1_RVT S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  FADDX1_RVT S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  FADDX1_RVT S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  FADDX1_RVT S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), 
        .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  FADDX1_RVT S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  FADDX1_RVT S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  FADDX1_RVT S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  FADDX1_RVT S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  FADDX1_RVT S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  FADDX1_RVT S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  FADDX1_RVT S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), 
        .S(SUMB_12__19_) );
  FADDX1_RVT S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(PRODUCT_11_) );
  FADDX1_RVT S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  FADDX1_RVT S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  FADDX1_RVT S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  FADDX1_RVT S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  FADDX1_RVT S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  FADDX1_RVT S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  FADDX1_RVT S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  FADDX1_RVT S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  FADDX1_RVT S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  FADDX1_RVT S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  FADDX1_RVT S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), 
        .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  FADDX1_RVT S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  FADDX1_RVT S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  FADDX1_RVT S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  FADDX1_RVT S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  FADDX1_RVT S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  FADDX1_RVT S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  FADDX1_RVT S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  FADDX1_RVT S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  FADDX1_RVT S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), 
        .S(SUMB_11__20_) );
  FADDX1_RVT S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT_10_) );
  FADDX1_RVT S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FADDX1_RVT S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FADDX1_RVT S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FADDX1_RVT S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FADDX1_RVT S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FADDX1_RVT S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FADDX1_RVT S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FADDX1_RVT S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FADDX1_RVT S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FADDX1_RVT S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  FADDX1_RVT S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  FADDX1_RVT S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  FADDX1_RVT S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  FADDX1_RVT S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  FADDX1_RVT S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  FADDX1_RVT S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  FADDX1_RVT S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  FADDX1_RVT S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  FADDX1_RVT S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  FADDX1_RVT S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  FADDX1_RVT S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .S(SUMB_10__21_) );
  FADDX1_RVT S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT_9_) );
  FADDX1_RVT S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FADDX1_RVT S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FADDX1_RVT S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FADDX1_RVT S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FADDX1_RVT S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FADDX1_RVT S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FADDX1_RVT S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FADDX1_RVT S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FADDX1_RVT S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FADDX1_RVT S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  FADDX1_RVT S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  FADDX1_RVT S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  FADDX1_RVT S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  FADDX1_RVT S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  FADDX1_RVT S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  FADDX1_RVT S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  FADDX1_RVT S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  FADDX1_RVT S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  FADDX1_RVT S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  FADDX1_RVT S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  FADDX1_RVT S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  FADDX1_RVT S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .S(
        SUMB_9__22_) );
  FADDX1_RVT S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT_8_) );
  FADDX1_RVT S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FADDX1_RVT S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FADDX1_RVT S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FADDX1_RVT S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FADDX1_RVT S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FADDX1_RVT S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FADDX1_RVT S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FADDX1_RVT S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FADDX1_RVT S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FADDX1_RVT S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  FADDX1_RVT S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  FADDX1_RVT S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  FADDX1_RVT S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  FADDX1_RVT S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  FADDX1_RVT S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  FADDX1_RVT S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  FADDX1_RVT S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  FADDX1_RVT S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  FADDX1_RVT S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  FADDX1_RVT S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  FADDX1_RVT S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  FADDX1_RVT S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  FADDX1_RVT S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .S(
        SUMB_8__23_) );
  FADDX1_RVT S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT_7_) );
  FADDX1_RVT S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FADDX1_RVT S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FADDX1_RVT S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FADDX1_RVT S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FADDX1_RVT S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FADDX1_RVT S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FADDX1_RVT S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FADDX1_RVT S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FADDX1_RVT S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FADDX1_RVT S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  FADDX1_RVT S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  FADDX1_RVT S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  FADDX1_RVT S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  FADDX1_RVT S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  FADDX1_RVT S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  FADDX1_RVT S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  FADDX1_RVT S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  FADDX1_RVT S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  FADDX1_RVT S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  FADDX1_RVT S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  FADDX1_RVT S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  FADDX1_RVT S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  FADDX1_RVT S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  FADDX1_RVT S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .S(
        SUMB_7__24_) );
  FADDX1_RVT S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT_6_) );
  FADDX1_RVT S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FADDX1_RVT S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FADDX1_RVT S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FADDX1_RVT S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FADDX1_RVT S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FADDX1_RVT S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FADDX1_RVT S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FADDX1_RVT S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FADDX1_RVT S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FADDX1_RVT S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  FADDX1_RVT S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  FADDX1_RVT S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  FADDX1_RVT S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  FADDX1_RVT S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  FADDX1_RVT S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  FADDX1_RVT S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  FADDX1_RVT S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  FADDX1_RVT S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  FADDX1_RVT S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  FADDX1_RVT S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  FADDX1_RVT S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  FADDX1_RVT S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  FADDX1_RVT S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  FADDX1_RVT S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  FADDX1_RVT S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .S(
        SUMB_6__25_) );
  FADDX1_RVT S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT_5_) );
  FADDX1_RVT S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FADDX1_RVT S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FADDX1_RVT S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FADDX1_RVT S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FADDX1_RVT S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FADDX1_RVT S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FADDX1_RVT S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FADDX1_RVT S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FADDX1_RVT S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FADDX1_RVT S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  FADDX1_RVT S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  FADDX1_RVT S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  FADDX1_RVT S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  FADDX1_RVT S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  FADDX1_RVT S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  FADDX1_RVT S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  FADDX1_RVT S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  FADDX1_RVT S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  FADDX1_RVT S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  FADDX1_RVT S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  FADDX1_RVT S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  FADDX1_RVT S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  FADDX1_RVT S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  FADDX1_RVT S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  FADDX1_RVT S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  FADDX1_RVT S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .S(
        SUMB_5__26_) );
  FADDX1_RVT S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT_4_) );
  FADDX1_RVT S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FADDX1_RVT S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FADDX1_RVT S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FADDX1_RVT S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FADDX1_RVT S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FADDX1_RVT S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FADDX1_RVT S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FADDX1_RVT S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FADDX1_RVT S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FADDX1_RVT S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  FADDX1_RVT S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  FADDX1_RVT S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  FADDX1_RVT S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  FADDX1_RVT S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  FADDX1_RVT S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  FADDX1_RVT S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  FADDX1_RVT S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  FADDX1_RVT S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  FADDX1_RVT S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  FADDX1_RVT S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  FADDX1_RVT S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  FADDX1_RVT S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  FADDX1_RVT S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  FADDX1_RVT S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  FADDX1_RVT S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  FADDX1_RVT S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  FADDX1_RVT S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .S(
        SUMB_4__27_) );
  FADDX1_RVT S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT_3_) );
  FADDX1_RVT S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FADDX1_RVT S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FADDX1_RVT S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FADDX1_RVT S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FADDX1_RVT S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FADDX1_RVT S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FADDX1_RVT S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FADDX1_RVT S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FADDX1_RVT S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FADDX1_RVT S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  FADDX1_RVT S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  FADDX1_RVT S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  FADDX1_RVT S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  FADDX1_RVT S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  FADDX1_RVT S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  FADDX1_RVT S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  FADDX1_RVT S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  FADDX1_RVT S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  FADDX1_RVT S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  FADDX1_RVT S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  FADDX1_RVT S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  FADDX1_RVT S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  FADDX1_RVT S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  FADDX1_RVT S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  FADDX1_RVT S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  FADDX1_RVT S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  FADDX1_RVT S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  FADDX1_RVT S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .S(
        SUMB_3__28_) );
  FADDX1_RVT S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(PRODUCT_2_) );
  FADDX1_RVT S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FADDX1_RVT S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FADDX1_RVT S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FADDX1_RVT S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FADDX1_RVT S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FADDX1_RVT S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FADDX1_RVT S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FADDX1_RVT S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FADDX1_RVT S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FADDX1_RVT S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), 
        .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  FADDX1_RVT S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), 
        .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  FADDX1_RVT S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), 
        .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  FADDX1_RVT S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), 
        .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  FADDX1_RVT S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), 
        .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  FADDX1_RVT S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), 
        .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  FADDX1_RVT S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), 
        .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  FADDX1_RVT S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), 
        .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  FADDX1_RVT S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), 
        .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  FADDX1_RVT S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), 
        .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  FADDX1_RVT S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), 
        .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  FADDX1_RVT S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), 
        .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  FADDX1_RVT S2_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(SUMB_1__23_), 
        .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  FADDX1_RVT S2_2_23 ( .A(ab_2__23_), .B(CARRYB_1__23_), .CI(SUMB_1__24_), 
        .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  FADDX1_RVT S2_2_24 ( .A(ab_2__24_), .B(CARRYB_1__24_), .CI(SUMB_1__25_), 
        .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  FADDX1_RVT S2_2_25 ( .A(ab_2__25_), .B(CARRYB_1__25_), .CI(SUMB_1__26_), 
        .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  FADDX1_RVT S2_2_26 ( .A(ab_2__26_), .B(CARRYB_1__26_), .CI(SUMB_1__27_), 
        .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  FADDX1_RVT S2_2_27 ( .A(ab_2__27_), .B(CARRYB_1__27_), .CI(SUMB_1__28_), 
        .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  FADDX1_RVT S2_2_28 ( .A(ab_2__28_), .B(CARRYB_1__28_), .CI(SUMB_1__29_), 
        .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  FADDX1_RVT S2_2_29 ( .A(ab_2__29_), .B(CARRYB_1__29_), .CI(SUMB_1__30_), .S(
        SUMB_2__29_) );
  XOR2X1_RVT U2 ( .A1(ab_0__3_), .A2(ab_1__2_), .Y(SUMB_1__2_) );
  XOR2X1_RVT U3 ( .A1(ab_0__6_), .A2(ab_1__5_), .Y(SUMB_1__5_) );
  XOR2X1_RVT U4 ( .A1(ab_0__5_), .A2(ab_1__4_), .Y(SUMB_1__4_) );
  XOR2X1_RVT U5 ( .A1(ab_0__4_), .A2(ab_1__3_), .Y(SUMB_1__3_) );
  XOR2X1_RVT U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .Y(SUMB_1__20_) );
  XOR2X1_RVT U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .Y(SUMB_1__19_) );
  XOR2X1_RVT U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .Y(SUMB_1__18_) );
  XOR2X1_RVT U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .Y(SUMB_1__17_) );
  XOR2X1_RVT U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .Y(SUMB_1__16_) );
  XOR2X1_RVT U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .Y(SUMB_1__15_) );
  XOR2X1_RVT U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .Y(SUMB_1__14_) );
  XOR2X1_RVT U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .Y(SUMB_1__13_) );
  XOR2X1_RVT U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .Y(SUMB_1__12_) );
  XOR2X1_RVT U15 ( .A1(ab_0__11_), .A2(ab_1__10_), .Y(SUMB_1__10_) );
  XOR2X1_RVT U16 ( .A1(ab_0__10_), .A2(ab_1__9_), .Y(SUMB_1__9_) );
  XOR2X1_RVT U17 ( .A1(ab_0__9_), .A2(ab_1__8_), .Y(SUMB_1__8_) );
  XOR2X1_RVT U18 ( .A1(ab_0__8_), .A2(ab_1__7_), .Y(SUMB_1__7_) );
  XOR2X1_RVT U19 ( .A1(ab_0__7_), .A2(ab_1__6_), .Y(SUMB_1__6_) );
  XOR2X1_RVT U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .Y(SUMB_1__21_) );
  XOR2X1_RVT U21 ( .A1(ab_0__2_), .A2(ab_1__1_), .Y(SUMB_1__1_) );
  XOR2X1_RVT U22 ( .A1(ab_0__12_), .A2(ab_1__11_), .Y(SUMB_1__11_) );
  NBUFFX2_RVT U23 ( .A(A[0]), .Y(n34) );
  NBUFFX2_RVT U24 ( .A(A[1]), .Y(n37) );
  NBUFFX2_RVT U25 ( .A(A[1]), .Y(n36) );
  NBUFFX2_RVT U26 ( .A(A[0]), .Y(n33) );
  NBUFFX2_RVT U27 ( .A(A[2]), .Y(n39) );
  NBUFFX2_RVT U28 ( .A(A[3]), .Y(n41) );
  XOR2X1_RVT U29 ( .A1(ab_0__31_), .A2(ab_1__30_), .Y(SUMB_1__30_) );
  NBUFFX2_RVT U30 ( .A(A[0]), .Y(n35) );
  NBUFFX2_RVT U31 ( .A(A[1]), .Y(n38) );
  XOR2X1_RVT U32 ( .A1(ab_0__30_), .A2(ab_1__29_), .Y(SUMB_1__29_) );
  XOR2X1_RVT U33 ( .A1(ab_0__29_), .A2(ab_1__28_), .Y(SUMB_1__28_) );
  XOR2X1_RVT U34 ( .A1(ab_0__28_), .A2(ab_1__27_), .Y(SUMB_1__27_) );
  XOR2X1_RVT U35 ( .A1(ab_0__27_), .A2(ab_1__26_), .Y(SUMB_1__26_) );
  XOR2X1_RVT U36 ( .A1(ab_0__26_), .A2(ab_1__25_), .Y(SUMB_1__25_) );
  XOR2X1_RVT U37 ( .A1(ab_0__25_), .A2(ab_1__24_), .Y(SUMB_1__24_) );
  XOR2X1_RVT U38 ( .A1(ab_0__24_), .A2(ab_1__23_), .Y(SUMB_1__23_) );
  XOR2X1_RVT U39 ( .A1(ab_0__23_), .A2(ab_1__22_), .Y(SUMB_1__22_) );
  NBUFFX2_RVT U40 ( .A(A[2]), .Y(n40) );
  NBUFFX2_RVT U41 ( .A(B[3]), .Y(n62) );
  NBUFFX2_RVT U42 ( .A(B[9]), .Y(n74) );
  NBUFFX2_RVT U43 ( .A(B[8]), .Y(n72) );
  NBUFFX2_RVT U44 ( .A(A[9]), .Y(n54) );
  NBUFFX2_RVT U45 ( .A(B[7]), .Y(n70) );
  NBUFFX2_RVT U46 ( .A(A[9]), .Y(n53) );
  NBUFFX2_RVT U47 ( .A(B[4]), .Y(n63) );
  NBUFFX2_RVT U48 ( .A(B[0]), .Y(n55) );
  NBUFFX2_RVT U49 ( .A(B[6]), .Y(n68) );
  NBUFFX2_RVT U50 ( .A(A[4]), .Y(n43) );
  NBUFFX2_RVT U51 ( .A(A[5]), .Y(n45) );
  NBUFFX2_RVT U52 ( .A(A[6]), .Y(n47) );
  NBUFFX2_RVT U53 ( .A(A[7]), .Y(n50) );
  NBUFFX2_RVT U54 ( .A(A[7]), .Y(n49) );
  NBUFFX2_RVT U55 ( .A(B[9]), .Y(n73) );
  NBUFFX2_RVT U56 ( .A(B[7]), .Y(n69) );
  NBUFFX2_RVT U57 ( .A(B[8]), .Y(n71) );
  NBUFFX2_RVT U58 ( .A(B[5]), .Y(n65) );
  NBUFFX2_RVT U59 ( .A(B[6]), .Y(n67) );
  NBUFFX2_RVT U60 ( .A(A[8]), .Y(n52) );
  NBUFFX2_RVT U61 ( .A(A[8]), .Y(n51) );
  NBUFFX2_RVT U62 ( .A(B[4]), .Y(n64) );
  NBUFFX2_RVT U63 ( .A(B[3]), .Y(n61) );
  NBUFFX2_RVT U64 ( .A(B[2]), .Y(n59) );
  NBUFFX2_RVT U65 ( .A(B[1]), .Y(n57) );
  NBUFFX2_RVT U66 ( .A(B[5]), .Y(n66) );
  XOR2X1_RVT U67 ( .A1(ab_0__1_), .A2(ab_1__0_), .Y(PRODUCT_1_) );
  NBUFFX2_RVT U68 ( .A(A[3]), .Y(n42) );
  NBUFFX2_RVT U69 ( .A(B[0]), .Y(n56) );
  NBUFFX2_RVT U70 ( .A(A[4]), .Y(n44) );
  NBUFFX2_RVT U71 ( .A(B[1]), .Y(n58) );
  NBUFFX2_RVT U72 ( .A(A[5]), .Y(n46) );
  NBUFFX2_RVT U73 ( .A(B[2]), .Y(n60) );
  NBUFFX2_RVT U74 ( .A(A[6]), .Y(n48) );
  AND2X1_RVT U75 ( .A1(ab_1__0_), .A2(ab_0__1_), .Y(CARRYB_1__0_) );
  AND2X1_RVT U76 ( .A1(ab_1__1_), .A2(ab_0__2_), .Y(CARRYB_1__1_) );
  AND2X1_RVT U77 ( .A1(ab_1__2_), .A2(ab_0__3_), .Y(CARRYB_1__2_) );
  AND2X1_RVT U78 ( .A1(ab_1__3_), .A2(ab_0__4_), .Y(CARRYB_1__3_) );
  AND2X1_RVT U79 ( .A1(ab_1__4_), .A2(ab_0__5_), .Y(CARRYB_1__4_) );
  AND2X1_RVT U80 ( .A1(ab_1__5_), .A2(ab_0__6_), .Y(CARRYB_1__5_) );
  AND2X1_RVT U81 ( .A1(ab_1__6_), .A2(ab_0__7_), .Y(CARRYB_1__6_) );
  AND2X1_RVT U82 ( .A1(ab_1__7_), .A2(ab_0__8_), .Y(CARRYB_1__7_) );
  AND2X1_RVT U83 ( .A1(ab_1__8_), .A2(ab_0__9_), .Y(CARRYB_1__8_) );
  AND2X1_RVT U84 ( .A1(ab_1__9_), .A2(ab_0__10_), .Y(CARRYB_1__9_) );
  AND2X1_RVT U85 ( .A1(ab_1__10_), .A2(ab_0__11_), .Y(CARRYB_1__10_) );
  AND2X1_RVT U86 ( .A1(ab_1__11_), .A2(ab_0__12_), .Y(CARRYB_1__11_) );
  AND2X1_RVT U87 ( .A1(ab_1__12_), .A2(ab_0__13_), .Y(CARRYB_1__12_) );
  AND2X1_RVT U88 ( .A1(ab_1__13_), .A2(ab_0__14_), .Y(CARRYB_1__13_) );
  AND2X1_RVT U89 ( .A1(ab_1__14_), .A2(ab_0__15_), .Y(CARRYB_1__14_) );
  AND2X1_RVT U90 ( .A1(ab_1__15_), .A2(ab_0__16_), .Y(CARRYB_1__15_) );
  AND2X1_RVT U91 ( .A1(ab_1__16_), .A2(ab_0__17_), .Y(CARRYB_1__16_) );
  AND2X1_RVT U92 ( .A1(ab_1__17_), .A2(ab_0__18_), .Y(CARRYB_1__17_) );
  AND2X1_RVT U93 ( .A1(ab_1__18_), .A2(ab_0__19_), .Y(CARRYB_1__18_) );
  AND2X1_RVT U94 ( .A1(ab_1__19_), .A2(ab_0__20_), .Y(CARRYB_1__19_) );
  AND2X1_RVT U95 ( .A1(ab_1__20_), .A2(ab_0__21_), .Y(CARRYB_1__20_) );
  AND2X1_RVT U96 ( .A1(ab_1__21_), .A2(ab_0__22_), .Y(CARRYB_1__21_) );
  AND2X1_RVT U97 ( .A1(ab_1__22_), .A2(ab_0__23_), .Y(CARRYB_1__22_) );
  AND2X1_RVT U98 ( .A1(ab_1__23_), .A2(ab_0__24_), .Y(CARRYB_1__23_) );
  AND2X1_RVT U99 ( .A1(ab_1__24_), .A2(ab_0__25_), .Y(CARRYB_1__24_) );
  AND2X1_RVT U100 ( .A1(ab_1__25_), .A2(ab_0__26_), .Y(CARRYB_1__25_) );
  AND2X1_RVT U101 ( .A1(ab_1__26_), .A2(ab_0__27_), .Y(CARRYB_1__26_) );
  AND2X1_RVT U102 ( .A1(ab_1__27_), .A2(ab_0__28_), .Y(CARRYB_1__27_) );
  AND2X1_RVT U103 ( .A1(ab_1__28_), .A2(ab_0__29_), .Y(CARRYB_1__28_) );
  AND2X1_RVT U104 ( .A1(ab_1__29_), .A2(ab_0__30_), .Y(CARRYB_1__29_) );
  NBUFFX2_RVT U105 ( .A(B[10]), .Y(n3) );
  NBUFFX2_RVT U106 ( .A(B[10]), .Y(n4) );
  NBUFFX2_RVT U107 ( .A(B[11]), .Y(n5) );
  NBUFFX2_RVT U108 ( .A(B[11]), .Y(n6) );
  NBUFFX2_RVT U109 ( .A(B[12]), .Y(n7) );
  NBUFFX2_RVT U110 ( .A(B[13]), .Y(n8) );
  NBUFFX2_RVT U111 ( .A(B[14]), .Y(n9) );
  NBUFFX2_RVT U112 ( .A(B[15]), .Y(n10) );
  NBUFFX2_RVT U113 ( .A(B[16]), .Y(n11) );
  NBUFFX2_RVT U114 ( .A(B[17]), .Y(n12) );
  NBUFFX2_RVT U115 ( .A(B[18]), .Y(n13) );
  INVX0_RVT U116 ( .A(B[19]), .Y(n14) );
  INVX0_RVT U117 ( .A(n14), .Y(n15) );
  INVX0_RVT U118 ( .A(B[20]), .Y(n16) );
  INVX0_RVT U119 ( .A(n16), .Y(n17) );
  NBUFFX2_RVT U120 ( .A(A[10]), .Y(n18) );
  NBUFFX2_RVT U121 ( .A(A[10]), .Y(n19) );
  NBUFFX2_RVT U122 ( .A(A[11]), .Y(n20) );
  NBUFFX2_RVT U123 ( .A(A[12]), .Y(n21) );
  NBUFFX2_RVT U124 ( .A(A[13]), .Y(n22) );
  NBUFFX2_RVT U125 ( .A(A[14]), .Y(n23) );
  NBUFFX2_RVT U126 ( .A(A[15]), .Y(n24) );
  NBUFFX2_RVT U127 ( .A(A[16]), .Y(n25) );
  NBUFFX2_RVT U128 ( .A(A[17]), .Y(n26) );
  NBUFFX2_RVT U129 ( .A(A[18]), .Y(n27) );
  NBUFFX2_RVT U130 ( .A(A[19]), .Y(n28) );
  INVX0_RVT U131 ( .A(A[20]), .Y(n29) );
  INVX0_RVT U132 ( .A(n29), .Y(n30) );
  INVX0_RVT U133 ( .A(A[21]), .Y(n31) );
  INVX0_RVT U134 ( .A(n31), .Y(n32) );
  AND2X1_RVT U135 ( .A1(n73), .A2(n54), .Y(ab_9__9_) );
  AND2X1_RVT U136 ( .A1(n71), .A2(n54), .Y(ab_9__8_) );
  AND2X1_RVT U137 ( .A1(n69), .A2(n54), .Y(ab_9__7_) );
  AND2X1_RVT U138 ( .A1(n67), .A2(n54), .Y(ab_9__6_) );
  AND2X1_RVT U139 ( .A1(n65), .A2(n54), .Y(ab_9__5_) );
  AND2X1_RVT U140 ( .A1(n63), .A2(n54), .Y(ab_9__4_) );
  AND2X1_RVT U141 ( .A1(n62), .A2(n54), .Y(ab_9__3_) );
  AND2X1_RVT U142 ( .A1(n60), .A2(n54), .Y(ab_9__2_) );
  AND2X1_RVT U143 ( .A1(B[22]), .A2(n54), .Y(ab_9__22_) );
  AND2X1_RVT U144 ( .A1(B[21]), .A2(n54), .Y(ab_9__21_) );
  AND2X1_RVT U145 ( .A1(n17), .A2(n54), .Y(ab_9__20_) );
  AND2X1_RVT U146 ( .A1(n58), .A2(n53), .Y(ab_9__1_) );
  AND2X1_RVT U147 ( .A1(n15), .A2(n53), .Y(ab_9__19_) );
  AND2X1_RVT U148 ( .A1(n13), .A2(n53), .Y(ab_9__18_) );
  AND2X1_RVT U149 ( .A1(B[17]), .A2(n53), .Y(ab_9__17_) );
  AND2X1_RVT U150 ( .A1(n11), .A2(n53), .Y(ab_9__16_) );
  AND2X1_RVT U151 ( .A1(n10), .A2(n53), .Y(ab_9__15_) );
  AND2X1_RVT U152 ( .A1(n9), .A2(n53), .Y(ab_9__14_) );
  AND2X1_RVT U153 ( .A1(B[13]), .A2(n53), .Y(ab_9__13_) );
  AND2X1_RVT U154 ( .A1(n7), .A2(n53), .Y(ab_9__12_) );
  AND2X1_RVT U155 ( .A1(n5), .A2(n53), .Y(ab_9__11_) );
  AND2X1_RVT U156 ( .A1(n3), .A2(n53), .Y(ab_9__10_) );
  AND2X1_RVT U157 ( .A1(n55), .A2(n53), .Y(ab_9__0_) );
  AND2X1_RVT U158 ( .A1(n52), .A2(n73), .Y(ab_8__9_) );
  AND2X1_RVT U159 ( .A1(n52), .A2(n71), .Y(ab_8__8_) );
  AND2X1_RVT U160 ( .A1(n52), .A2(n69), .Y(ab_8__7_) );
  AND2X1_RVT U161 ( .A1(n52), .A2(n67), .Y(ab_8__6_) );
  AND2X1_RVT U162 ( .A1(n52), .A2(n65), .Y(ab_8__5_) );
  AND2X1_RVT U163 ( .A1(n52), .A2(n63), .Y(ab_8__4_) );
  AND2X1_RVT U164 ( .A1(n52), .A2(n62), .Y(ab_8__3_) );
  AND2X1_RVT U165 ( .A1(n52), .A2(n60), .Y(ab_8__2_) );
  AND2X1_RVT U166 ( .A1(n52), .A2(B[23]), .Y(ab_8__23_) );
  AND2X1_RVT U167 ( .A1(n52), .A2(B[22]), .Y(ab_8__22_) );
  AND2X1_RVT U168 ( .A1(n52), .A2(B[21]), .Y(ab_8__21_) );
  AND2X1_RVT U169 ( .A1(n52), .A2(n17), .Y(ab_8__20_) );
  AND2X1_RVT U170 ( .A1(n51), .A2(n58), .Y(ab_8__1_) );
  AND2X1_RVT U171 ( .A1(n51), .A2(n15), .Y(ab_8__19_) );
  AND2X1_RVT U172 ( .A1(n51), .A2(n13), .Y(ab_8__18_) );
  AND2X1_RVT U173 ( .A1(n51), .A2(n12), .Y(ab_8__17_) );
  AND2X1_RVT U174 ( .A1(n51), .A2(n11), .Y(ab_8__16_) );
  AND2X1_RVT U175 ( .A1(n51), .A2(n10), .Y(ab_8__15_) );
  AND2X1_RVT U176 ( .A1(n51), .A2(n9), .Y(ab_8__14_) );
  AND2X1_RVT U177 ( .A1(n51), .A2(B[13]), .Y(ab_8__13_) );
  AND2X1_RVT U178 ( .A1(n51), .A2(n7), .Y(ab_8__12_) );
  AND2X1_RVT U179 ( .A1(n51), .A2(n5), .Y(ab_8__11_) );
  AND2X1_RVT U180 ( .A1(n51), .A2(n4), .Y(ab_8__10_) );
  AND2X1_RVT U181 ( .A1(n51), .A2(n55), .Y(ab_8__0_) );
  AND2X1_RVT U182 ( .A1(n49), .A2(n73), .Y(ab_7__9_) );
  AND2X1_RVT U183 ( .A1(n50), .A2(n71), .Y(ab_7__8_) );
  AND2X1_RVT U184 ( .A1(n50), .A2(n69), .Y(ab_7__7_) );
  AND2X1_RVT U185 ( .A1(n50), .A2(n67), .Y(ab_7__6_) );
  AND2X1_RVT U186 ( .A1(n50), .A2(n65), .Y(ab_7__5_) );
  AND2X1_RVT U187 ( .A1(n50), .A2(n63), .Y(ab_7__4_) );
  AND2X1_RVT U188 ( .A1(n50), .A2(n62), .Y(ab_7__3_) );
  AND2X1_RVT U189 ( .A1(n50), .A2(n60), .Y(ab_7__2_) );
  AND2X1_RVT U190 ( .A1(n50), .A2(B[24]), .Y(ab_7__24_) );
  AND2X1_RVT U191 ( .A1(n50), .A2(B[23]), .Y(ab_7__23_) );
  AND2X1_RVT U192 ( .A1(n50), .A2(B[22]), .Y(ab_7__22_) );
  AND2X1_RVT U193 ( .A1(n50), .A2(B[21]), .Y(ab_7__21_) );
  AND2X1_RVT U194 ( .A1(n50), .A2(n17), .Y(ab_7__20_) );
  AND2X1_RVT U195 ( .A1(n49), .A2(n58), .Y(ab_7__1_) );
  AND2X1_RVT U196 ( .A1(n49), .A2(n15), .Y(ab_7__19_) );
  AND2X1_RVT U197 ( .A1(n49), .A2(n13), .Y(ab_7__18_) );
  AND2X1_RVT U198 ( .A1(n49), .A2(n12), .Y(ab_7__17_) );
  AND2X1_RVT U199 ( .A1(n49), .A2(n11), .Y(ab_7__16_) );
  AND2X1_RVT U200 ( .A1(n49), .A2(n10), .Y(ab_7__15_) );
  AND2X1_RVT U201 ( .A1(n49), .A2(n9), .Y(ab_7__14_) );
  AND2X1_RVT U202 ( .A1(n49), .A2(B[13]), .Y(ab_7__13_) );
  AND2X1_RVT U203 ( .A1(n49), .A2(n7), .Y(ab_7__12_) );
  AND2X1_RVT U204 ( .A1(n49), .A2(n5), .Y(ab_7__11_) );
  AND2X1_RVT U205 ( .A1(n49), .A2(n3), .Y(ab_7__10_) );
  AND2X1_RVT U206 ( .A1(n49), .A2(n55), .Y(ab_7__0_) );
  AND2X1_RVT U207 ( .A1(n48), .A2(n73), .Y(ab_6__9_) );
  AND2X1_RVT U208 ( .A1(n48), .A2(n71), .Y(ab_6__8_) );
  AND2X1_RVT U209 ( .A1(n47), .A2(n69), .Y(ab_6__7_) );
  AND2X1_RVT U210 ( .A1(n47), .A2(n67), .Y(ab_6__6_) );
  AND2X1_RVT U211 ( .A1(n47), .A2(n65), .Y(ab_6__5_) );
  AND2X1_RVT U212 ( .A1(n47), .A2(n63), .Y(ab_6__4_) );
  AND2X1_RVT U213 ( .A1(n47), .A2(n62), .Y(ab_6__3_) );
  AND2X1_RVT U214 ( .A1(n47), .A2(n60), .Y(ab_6__2_) );
  AND2X1_RVT U215 ( .A1(n47), .A2(B[25]), .Y(ab_6__25_) );
  AND2X1_RVT U216 ( .A1(n47), .A2(B[24]), .Y(ab_6__24_) );
  AND2X1_RVT U217 ( .A1(n47), .A2(B[23]), .Y(ab_6__23_) );
  AND2X1_RVT U218 ( .A1(n47), .A2(B[22]), .Y(ab_6__22_) );
  AND2X1_RVT U219 ( .A1(n47), .A2(B[21]), .Y(ab_6__21_) );
  AND2X1_RVT U220 ( .A1(n47), .A2(n17), .Y(ab_6__20_) );
  AND2X1_RVT U221 ( .A1(n48), .A2(n58), .Y(ab_6__1_) );
  AND2X1_RVT U222 ( .A1(n48), .A2(n15), .Y(ab_6__19_) );
  AND2X1_RVT U223 ( .A1(n48), .A2(n13), .Y(ab_6__18_) );
  AND2X1_RVT U224 ( .A1(n48), .A2(n12), .Y(ab_6__17_) );
  AND2X1_RVT U225 ( .A1(n48), .A2(n11), .Y(ab_6__16_) );
  AND2X1_RVT U226 ( .A1(n48), .A2(n10), .Y(ab_6__15_) );
  AND2X1_RVT U227 ( .A1(n48), .A2(n9), .Y(ab_6__14_) );
  AND2X1_RVT U228 ( .A1(n48), .A2(n8), .Y(ab_6__13_) );
  AND2X1_RVT U229 ( .A1(n48), .A2(n7), .Y(ab_6__12_) );
  AND2X1_RVT U230 ( .A1(n48), .A2(n5), .Y(ab_6__11_) );
  AND2X1_RVT U231 ( .A1(n48), .A2(n4), .Y(ab_6__10_) );
  AND2X1_RVT U232 ( .A1(n48), .A2(n55), .Y(ab_6__0_) );
  AND2X1_RVT U233 ( .A1(n46), .A2(n73), .Y(ab_5__9_) );
  AND2X1_RVT U234 ( .A1(n46), .A2(n71), .Y(ab_5__8_) );
  AND2X1_RVT U235 ( .A1(n46), .A2(n69), .Y(ab_5__7_) );
  AND2X1_RVT U236 ( .A1(n45), .A2(n67), .Y(ab_5__6_) );
  AND2X1_RVT U237 ( .A1(n45), .A2(n65), .Y(ab_5__5_) );
  AND2X1_RVT U238 ( .A1(n45), .A2(n63), .Y(ab_5__4_) );
  AND2X1_RVT U239 ( .A1(n45), .A2(n62), .Y(ab_5__3_) );
  AND2X1_RVT U240 ( .A1(n45), .A2(n60), .Y(ab_5__2_) );
  AND2X1_RVT U241 ( .A1(n45), .A2(B[26]), .Y(ab_5__26_) );
  AND2X1_RVT U242 ( .A1(n45), .A2(B[25]), .Y(ab_5__25_) );
  AND2X1_RVT U243 ( .A1(n45), .A2(B[24]), .Y(ab_5__24_) );
  AND2X1_RVT U244 ( .A1(n45), .A2(B[23]), .Y(ab_5__23_) );
  AND2X1_RVT U245 ( .A1(n45), .A2(B[22]), .Y(ab_5__22_) );
  AND2X1_RVT U246 ( .A1(n45), .A2(B[21]), .Y(ab_5__21_) );
  AND2X1_RVT U247 ( .A1(n45), .A2(n17), .Y(ab_5__20_) );
  AND2X1_RVT U248 ( .A1(n46), .A2(n58), .Y(ab_5__1_) );
  AND2X1_RVT U249 ( .A1(n46), .A2(n15), .Y(ab_5__19_) );
  AND2X1_RVT U250 ( .A1(n46), .A2(n13), .Y(ab_5__18_) );
  AND2X1_RVT U251 ( .A1(n46), .A2(n12), .Y(ab_5__17_) );
  AND2X1_RVT U252 ( .A1(n46), .A2(n11), .Y(ab_5__16_) );
  AND2X1_RVT U253 ( .A1(n46), .A2(n10), .Y(ab_5__15_) );
  AND2X1_RVT U254 ( .A1(n46), .A2(n9), .Y(ab_5__14_) );
  AND2X1_RVT U255 ( .A1(n46), .A2(n8), .Y(ab_5__13_) );
  AND2X1_RVT U256 ( .A1(n46), .A2(n7), .Y(ab_5__12_) );
  AND2X1_RVT U257 ( .A1(n46), .A2(n5), .Y(ab_5__11_) );
  AND2X1_RVT U258 ( .A1(n46), .A2(n3), .Y(ab_5__10_) );
  AND2X1_RVT U259 ( .A1(n46), .A2(n55), .Y(ab_5__0_) );
  AND2X1_RVT U260 ( .A1(n44), .A2(n73), .Y(ab_4__9_) );
  AND2X1_RVT U261 ( .A1(n44), .A2(n71), .Y(ab_4__8_) );
  AND2X1_RVT U262 ( .A1(n44), .A2(n69), .Y(ab_4__7_) );
  AND2X1_RVT U263 ( .A1(n44), .A2(n67), .Y(ab_4__6_) );
  AND2X1_RVT U264 ( .A1(n43), .A2(n65), .Y(ab_4__5_) );
  AND2X1_RVT U265 ( .A1(n43), .A2(n63), .Y(ab_4__4_) );
  AND2X1_RVT U266 ( .A1(n43), .A2(n62), .Y(ab_4__3_) );
  AND2X1_RVT U267 ( .A1(n43), .A2(n60), .Y(ab_4__2_) );
  AND2X1_RVT U268 ( .A1(n43), .A2(B[27]), .Y(ab_4__27_) );
  AND2X1_RVT U269 ( .A1(n43), .A2(B[26]), .Y(ab_4__26_) );
  AND2X1_RVT U270 ( .A1(n43), .A2(B[25]), .Y(ab_4__25_) );
  AND2X1_RVT U271 ( .A1(n43), .A2(B[24]), .Y(ab_4__24_) );
  AND2X1_RVT U272 ( .A1(n43), .A2(B[23]), .Y(ab_4__23_) );
  AND2X1_RVT U273 ( .A1(n43), .A2(B[22]), .Y(ab_4__22_) );
  AND2X1_RVT U274 ( .A1(n43), .A2(B[21]), .Y(ab_4__21_) );
  AND2X1_RVT U275 ( .A1(n43), .A2(n17), .Y(ab_4__20_) );
  AND2X1_RVT U276 ( .A1(n44), .A2(n58), .Y(ab_4__1_) );
  AND2X1_RVT U277 ( .A1(n44), .A2(n15), .Y(ab_4__19_) );
  AND2X1_RVT U278 ( .A1(n44), .A2(n13), .Y(ab_4__18_) );
  AND2X1_RVT U279 ( .A1(n44), .A2(n12), .Y(ab_4__17_) );
  AND2X1_RVT U280 ( .A1(n44), .A2(n11), .Y(ab_4__16_) );
  AND2X1_RVT U281 ( .A1(n44), .A2(n10), .Y(ab_4__15_) );
  AND2X1_RVT U282 ( .A1(n44), .A2(n9), .Y(ab_4__14_) );
  AND2X1_RVT U283 ( .A1(n44), .A2(n8), .Y(ab_4__13_) );
  AND2X1_RVT U284 ( .A1(n44), .A2(n7), .Y(ab_4__12_) );
  AND2X1_RVT U285 ( .A1(n44), .A2(n5), .Y(ab_4__11_) );
  AND2X1_RVT U286 ( .A1(n44), .A2(n4), .Y(ab_4__10_) );
  AND2X1_RVT U287 ( .A1(n44), .A2(n55), .Y(ab_4__0_) );
  AND2X1_RVT U288 ( .A1(n42), .A2(n73), .Y(ab_3__9_) );
  AND2X1_RVT U289 ( .A1(n42), .A2(n71), .Y(ab_3__8_) );
  AND2X1_RVT U290 ( .A1(n42), .A2(n69), .Y(ab_3__7_) );
  AND2X1_RVT U291 ( .A1(n42), .A2(n67), .Y(ab_3__6_) );
  AND2X1_RVT U292 ( .A1(n42), .A2(n65), .Y(ab_3__5_) );
  AND2X1_RVT U293 ( .A1(n41), .A2(n63), .Y(ab_3__4_) );
  AND2X1_RVT U294 ( .A1(n41), .A2(n62), .Y(ab_3__3_) );
  AND2X1_RVT U295 ( .A1(n41), .A2(n60), .Y(ab_3__2_) );
  AND2X1_RVT U296 ( .A1(n41), .A2(B[28]), .Y(ab_3__28_) );
  AND2X1_RVT U297 ( .A1(n41), .A2(B[27]), .Y(ab_3__27_) );
  AND2X1_RVT U298 ( .A1(n41), .A2(B[26]), .Y(ab_3__26_) );
  AND2X1_RVT U299 ( .A1(n41), .A2(B[25]), .Y(ab_3__25_) );
  AND2X1_RVT U300 ( .A1(n41), .A2(B[24]), .Y(ab_3__24_) );
  AND2X1_RVT U301 ( .A1(n41), .A2(B[23]), .Y(ab_3__23_) );
  AND2X1_RVT U302 ( .A1(n41), .A2(B[22]), .Y(ab_3__22_) );
  AND2X1_RVT U303 ( .A1(n41), .A2(B[21]), .Y(ab_3__21_) );
  AND2X1_RVT U304 ( .A1(n41), .A2(n17), .Y(ab_3__20_) );
  AND2X1_RVT U305 ( .A1(n42), .A2(n58), .Y(ab_3__1_) );
  AND2X1_RVT U306 ( .A1(n42), .A2(n15), .Y(ab_3__19_) );
  AND2X1_RVT U307 ( .A1(n42), .A2(n13), .Y(ab_3__18_) );
  AND2X1_RVT U308 ( .A1(n42), .A2(n12), .Y(ab_3__17_) );
  AND2X1_RVT U309 ( .A1(n42), .A2(n11), .Y(ab_3__16_) );
  AND2X1_RVT U310 ( .A1(n42), .A2(n10), .Y(ab_3__15_) );
  AND2X1_RVT U311 ( .A1(n42), .A2(n9), .Y(ab_3__14_) );
  AND2X1_RVT U312 ( .A1(n42), .A2(n8), .Y(ab_3__13_) );
  AND2X1_RVT U313 ( .A1(n42), .A2(n7), .Y(ab_3__12_) );
  AND2X1_RVT U314 ( .A1(n42), .A2(n5), .Y(ab_3__11_) );
  AND2X1_RVT U315 ( .A1(n42), .A2(n3), .Y(ab_3__10_) );
  AND2X1_RVT U316 ( .A1(n42), .A2(n55), .Y(ab_3__0_) );
  AND2X1_RVT U317 ( .A1(A[31]), .A2(n55), .Y(ab_31__0_) );
  AND2X1_RVT U318 ( .A1(A[30]), .A2(n58), .Y(ab_30__1_) );
  AND2X1_RVT U319 ( .A1(A[30]), .A2(n55), .Y(ab_30__0_) );
  AND2X1_RVT U320 ( .A1(n40), .A2(n73), .Y(ab_2__9_) );
  AND2X1_RVT U321 ( .A1(n40), .A2(n71), .Y(ab_2__8_) );
  AND2X1_RVT U322 ( .A1(n40), .A2(n69), .Y(ab_2__7_) );
  AND2X1_RVT U323 ( .A1(n40), .A2(n67), .Y(ab_2__6_) );
  AND2X1_RVT U324 ( .A1(n40), .A2(n65), .Y(ab_2__5_) );
  AND2X1_RVT U325 ( .A1(n40), .A2(n63), .Y(ab_2__4_) );
  AND2X1_RVT U326 ( .A1(n40), .A2(n62), .Y(ab_2__3_) );
  AND2X1_RVT U327 ( .A1(A[2]), .A2(n60), .Y(ab_2__2_) );
  AND2X1_RVT U328 ( .A1(A[2]), .A2(B[29]), .Y(ab_2__29_) );
  AND2X1_RVT U329 ( .A1(A[2]), .A2(B[28]), .Y(ab_2__28_) );
  AND2X1_RVT U330 ( .A1(n40), .A2(B[27]), .Y(ab_2__27_) );
  AND2X1_RVT U331 ( .A1(n39), .A2(B[26]), .Y(ab_2__26_) );
  AND2X1_RVT U332 ( .A1(n39), .A2(B[25]), .Y(ab_2__25_) );
  AND2X1_RVT U333 ( .A1(A[2]), .A2(B[24]), .Y(ab_2__24_) );
  AND2X1_RVT U334 ( .A1(n40), .A2(B[23]), .Y(ab_2__23_) );
  AND2X1_RVT U335 ( .A1(n39), .A2(B[22]), .Y(ab_2__22_) );
  AND2X1_RVT U336 ( .A1(A[2]), .A2(B[21]), .Y(ab_2__21_) );
  AND2X1_RVT U337 ( .A1(A[2]), .A2(n17), .Y(ab_2__20_) );
  AND2X1_RVT U338 ( .A1(n39), .A2(n58), .Y(ab_2__1_) );
  AND2X1_RVT U339 ( .A1(n39), .A2(n15), .Y(ab_2__19_) );
  AND2X1_RVT U340 ( .A1(n39), .A2(n13), .Y(ab_2__18_) );
  AND2X1_RVT U341 ( .A1(n39), .A2(n12), .Y(ab_2__17_) );
  AND2X1_RVT U342 ( .A1(n39), .A2(n11), .Y(ab_2__16_) );
  AND2X1_RVT U343 ( .A1(n39), .A2(n10), .Y(ab_2__15_) );
  AND2X1_RVT U344 ( .A1(n39), .A2(n9), .Y(ab_2__14_) );
  AND2X1_RVT U345 ( .A1(n39), .A2(n8), .Y(ab_2__13_) );
  AND2X1_RVT U346 ( .A1(n39), .A2(n7), .Y(ab_2__12_) );
  AND2X1_RVT U347 ( .A1(n39), .A2(n5), .Y(ab_2__11_) );
  AND2X1_RVT U348 ( .A1(n39), .A2(n4), .Y(ab_2__10_) );
  AND2X1_RVT U349 ( .A1(n39), .A2(n55), .Y(ab_2__0_) );
  AND2X1_RVT U350 ( .A1(A[29]), .A2(n60), .Y(ab_29__2_) );
  AND2X1_RVT U351 ( .A1(A[29]), .A2(n58), .Y(ab_29__1_) );
  AND2X1_RVT U352 ( .A1(A[29]), .A2(n55), .Y(ab_29__0_) );
  AND2X1_RVT U353 ( .A1(A[28]), .A2(n62), .Y(ab_28__3_) );
  AND2X1_RVT U354 ( .A1(A[28]), .A2(n60), .Y(ab_28__2_) );
  AND2X1_RVT U355 ( .A1(A[28]), .A2(n58), .Y(ab_28__1_) );
  AND2X1_RVT U356 ( .A1(A[28]), .A2(n55), .Y(ab_28__0_) );
  AND2X1_RVT U357 ( .A1(A[27]), .A2(n63), .Y(ab_27__4_) );
  AND2X1_RVT U358 ( .A1(A[27]), .A2(n62), .Y(ab_27__3_) );
  AND2X1_RVT U359 ( .A1(A[27]), .A2(n60), .Y(ab_27__2_) );
  AND2X1_RVT U360 ( .A1(A[27]), .A2(n58), .Y(ab_27__1_) );
  AND2X1_RVT U361 ( .A1(A[27]), .A2(n55), .Y(ab_27__0_) );
  AND2X1_RVT U362 ( .A1(A[26]), .A2(n65), .Y(ab_26__5_) );
  AND2X1_RVT U363 ( .A1(A[26]), .A2(n63), .Y(ab_26__4_) );
  AND2X1_RVT U364 ( .A1(A[26]), .A2(n62), .Y(ab_26__3_) );
  AND2X1_RVT U365 ( .A1(A[26]), .A2(n60), .Y(ab_26__2_) );
  AND2X1_RVT U366 ( .A1(A[26]), .A2(n58), .Y(ab_26__1_) );
  AND2X1_RVT U367 ( .A1(A[26]), .A2(n56), .Y(ab_26__0_) );
  AND2X1_RVT U368 ( .A1(A[25]), .A2(n67), .Y(ab_25__6_) );
  AND2X1_RVT U369 ( .A1(A[25]), .A2(n65), .Y(ab_25__5_) );
  AND2X1_RVT U370 ( .A1(A[25]), .A2(n63), .Y(ab_25__4_) );
  AND2X1_RVT U371 ( .A1(A[25]), .A2(n62), .Y(ab_25__3_) );
  AND2X1_RVT U372 ( .A1(A[25]), .A2(n60), .Y(ab_25__2_) );
  AND2X1_RVT U373 ( .A1(A[25]), .A2(n57), .Y(ab_25__1_) );
  AND2X1_RVT U374 ( .A1(A[25]), .A2(n56), .Y(ab_25__0_) );
  AND2X1_RVT U375 ( .A1(A[24]), .A2(n69), .Y(ab_24__7_) );
  AND2X1_RVT U376 ( .A1(A[24]), .A2(n67), .Y(ab_24__6_) );
  AND2X1_RVT U377 ( .A1(A[24]), .A2(n65), .Y(ab_24__5_) );
  AND2X1_RVT U378 ( .A1(A[24]), .A2(n63), .Y(ab_24__4_) );
  AND2X1_RVT U379 ( .A1(A[24]), .A2(n62), .Y(ab_24__3_) );
  AND2X1_RVT U380 ( .A1(A[24]), .A2(n59), .Y(ab_24__2_) );
  AND2X1_RVT U381 ( .A1(A[24]), .A2(n57), .Y(ab_24__1_) );
  AND2X1_RVT U382 ( .A1(A[24]), .A2(n56), .Y(ab_24__0_) );
  AND2X1_RVT U383 ( .A1(A[23]), .A2(n71), .Y(ab_23__8_) );
  AND2X1_RVT U384 ( .A1(A[23]), .A2(n69), .Y(ab_23__7_) );
  AND2X1_RVT U385 ( .A1(A[23]), .A2(n67), .Y(ab_23__6_) );
  AND2X1_RVT U386 ( .A1(A[23]), .A2(n65), .Y(ab_23__5_) );
  AND2X1_RVT U387 ( .A1(A[23]), .A2(n63), .Y(ab_23__4_) );
  AND2X1_RVT U388 ( .A1(A[23]), .A2(n61), .Y(ab_23__3_) );
  AND2X1_RVT U389 ( .A1(A[23]), .A2(n59), .Y(ab_23__2_) );
  AND2X1_RVT U390 ( .A1(A[23]), .A2(n57), .Y(ab_23__1_) );
  AND2X1_RVT U391 ( .A1(A[23]), .A2(n56), .Y(ab_23__0_) );
  AND2X1_RVT U392 ( .A1(A[22]), .A2(n73), .Y(ab_22__9_) );
  AND2X1_RVT U393 ( .A1(A[22]), .A2(n71), .Y(ab_22__8_) );
  AND2X1_RVT U394 ( .A1(A[22]), .A2(n69), .Y(ab_22__7_) );
  AND2X1_RVT U395 ( .A1(A[22]), .A2(n67), .Y(ab_22__6_) );
  AND2X1_RVT U396 ( .A1(A[22]), .A2(n65), .Y(ab_22__5_) );
  AND2X1_RVT U397 ( .A1(A[22]), .A2(n64), .Y(ab_22__4_) );
  AND2X1_RVT U398 ( .A1(A[22]), .A2(n61), .Y(ab_22__3_) );
  AND2X1_RVT U399 ( .A1(A[22]), .A2(n59), .Y(ab_22__2_) );
  AND2X1_RVT U400 ( .A1(A[22]), .A2(n57), .Y(ab_22__1_) );
  AND2X1_RVT U401 ( .A1(A[22]), .A2(n56), .Y(ab_22__0_) );
  AND2X1_RVT U402 ( .A1(A[21]), .A2(n73), .Y(ab_21__9_) );
  AND2X1_RVT U403 ( .A1(n32), .A2(n71), .Y(ab_21__8_) );
  AND2X1_RVT U404 ( .A1(n32), .A2(n69), .Y(ab_21__7_) );
  AND2X1_RVT U405 ( .A1(n32), .A2(n67), .Y(ab_21__6_) );
  AND2X1_RVT U406 ( .A1(n32), .A2(n66), .Y(ab_21__5_) );
  AND2X1_RVT U407 ( .A1(n32), .A2(n64), .Y(ab_21__4_) );
  AND2X1_RVT U408 ( .A1(n32), .A2(n61), .Y(ab_21__3_) );
  AND2X1_RVT U409 ( .A1(n32), .A2(n59), .Y(ab_21__2_) );
  AND2X1_RVT U410 ( .A1(n32), .A2(n57), .Y(ab_21__1_) );
  AND2X1_RVT U411 ( .A1(A[21]), .A2(n3), .Y(ab_21__10_) );
  AND2X1_RVT U412 ( .A1(n32), .A2(n56), .Y(ab_21__0_) );
  AND2X1_RVT U413 ( .A1(n30), .A2(n73), .Y(ab_20__9_) );
  AND2X1_RVT U414 ( .A1(n30), .A2(n71), .Y(ab_20__8_) );
  AND2X1_RVT U415 ( .A1(n30), .A2(n69), .Y(ab_20__7_) );
  AND2X1_RVT U416 ( .A1(n30), .A2(n68), .Y(ab_20__6_) );
  AND2X1_RVT U417 ( .A1(n30), .A2(n66), .Y(ab_20__5_) );
  AND2X1_RVT U418 ( .A1(n30), .A2(n64), .Y(ab_20__4_) );
  AND2X1_RVT U419 ( .A1(n30), .A2(n61), .Y(ab_20__3_) );
  AND2X1_RVT U420 ( .A1(n30), .A2(n59), .Y(ab_20__2_) );
  AND2X1_RVT U421 ( .A1(n30), .A2(n57), .Y(ab_20__1_) );
  AND2X1_RVT U422 ( .A1(A[20]), .A2(n5), .Y(ab_20__11_) );
  AND2X1_RVT U423 ( .A1(n30), .A2(n4), .Y(ab_20__10_) );
  AND2X1_RVT U424 ( .A1(n30), .A2(n56), .Y(ab_20__0_) );
  AND2X1_RVT U425 ( .A1(n38), .A2(n73), .Y(ab_1__9_) );
  AND2X1_RVT U426 ( .A1(n38), .A2(n71), .Y(ab_1__8_) );
  AND2X1_RVT U427 ( .A1(n38), .A2(n70), .Y(ab_1__7_) );
  AND2X1_RVT U428 ( .A1(n38), .A2(n68), .Y(ab_1__6_) );
  AND2X1_RVT U429 ( .A1(n38), .A2(n66), .Y(ab_1__5_) );
  AND2X1_RVT U430 ( .A1(n38), .A2(n64), .Y(ab_1__4_) );
  AND2X1_RVT U431 ( .A1(n38), .A2(n61), .Y(ab_1__3_) );
  AND2X1_RVT U432 ( .A1(n37), .A2(B[30]), .Y(ab_1__30_) );
  AND2X1_RVT U433 ( .A1(n37), .A2(n59), .Y(ab_1__2_) );
  AND2X1_RVT U434 ( .A1(n37), .A2(B[29]), .Y(ab_1__29_) );
  AND2X1_RVT U435 ( .A1(n37), .A2(B[28]), .Y(ab_1__28_) );
  AND2X1_RVT U436 ( .A1(n37), .A2(B[27]), .Y(ab_1__27_) );
  AND2X1_RVT U437 ( .A1(n37), .A2(B[26]), .Y(ab_1__26_) );
  AND2X1_RVT U438 ( .A1(n37), .A2(B[25]), .Y(ab_1__25_) );
  AND2X1_RVT U439 ( .A1(n37), .A2(B[24]), .Y(ab_1__24_) );
  AND2X1_RVT U440 ( .A1(n37), .A2(B[23]), .Y(ab_1__23_) );
  AND2X1_RVT U441 ( .A1(n37), .A2(B[22]), .Y(ab_1__22_) );
  AND2X1_RVT U442 ( .A1(n37), .A2(B[21]), .Y(ab_1__21_) );
  AND2X1_RVT U443 ( .A1(n37), .A2(B[20]), .Y(ab_1__20_) );
  AND2X1_RVT U444 ( .A1(n36), .A2(n57), .Y(ab_1__1_) );
  AND2X1_RVT U445 ( .A1(n36), .A2(B[19]), .Y(ab_1__19_) );
  AND2X1_RVT U446 ( .A1(n36), .A2(B[18]), .Y(ab_1__18_) );
  AND2X1_RVT U447 ( .A1(n36), .A2(n12), .Y(ab_1__17_) );
  AND2X1_RVT U448 ( .A1(n36), .A2(B[16]), .Y(ab_1__16_) );
  AND2X1_RVT U449 ( .A1(n36), .A2(B[15]), .Y(ab_1__15_) );
  AND2X1_RVT U450 ( .A1(n36), .A2(n9), .Y(ab_1__14_) );
  AND2X1_RVT U451 ( .A1(n36), .A2(B[13]), .Y(ab_1__13_) );
  AND2X1_RVT U452 ( .A1(n36), .A2(n7), .Y(ab_1__12_) );
  AND2X1_RVT U453 ( .A1(n36), .A2(n5), .Y(ab_1__11_) );
  AND2X1_RVT U454 ( .A1(n36), .A2(n3), .Y(ab_1__10_) );
  AND2X1_RVT U455 ( .A1(n36), .A2(B[0]), .Y(ab_1__0_) );
  AND2X1_RVT U456 ( .A1(n28), .A2(n73), .Y(ab_19__9_) );
  AND2X1_RVT U457 ( .A1(n28), .A2(n72), .Y(ab_19__8_) );
  AND2X1_RVT U458 ( .A1(n28), .A2(n70), .Y(ab_19__7_) );
  AND2X1_RVT U459 ( .A1(n28), .A2(n68), .Y(ab_19__6_) );
  AND2X1_RVT U460 ( .A1(n28), .A2(n66), .Y(ab_19__5_) );
  AND2X1_RVT U461 ( .A1(n28), .A2(n64), .Y(ab_19__4_) );
  AND2X1_RVT U462 ( .A1(n28), .A2(n61), .Y(ab_19__3_) );
  AND2X1_RVT U463 ( .A1(n28), .A2(n59), .Y(ab_19__2_) );
  AND2X1_RVT U464 ( .A1(n28), .A2(n57), .Y(ab_19__1_) );
  AND2X1_RVT U465 ( .A1(n28), .A2(B[12]), .Y(ab_19__12_) );
  AND2X1_RVT U466 ( .A1(n28), .A2(n6), .Y(ab_19__11_) );
  AND2X1_RVT U467 ( .A1(n28), .A2(n4), .Y(ab_19__10_) );
  AND2X1_RVT U468 ( .A1(A[19]), .A2(n56), .Y(ab_19__0_) );
  AND2X1_RVT U469 ( .A1(n27), .A2(n74), .Y(ab_18__9_) );
  AND2X1_RVT U470 ( .A1(n27), .A2(n72), .Y(ab_18__8_) );
  AND2X1_RVT U471 ( .A1(n27), .A2(n70), .Y(ab_18__7_) );
  AND2X1_RVT U472 ( .A1(n27), .A2(n68), .Y(ab_18__6_) );
  AND2X1_RVT U473 ( .A1(n27), .A2(n66), .Y(ab_18__5_) );
  AND2X1_RVT U474 ( .A1(n27), .A2(n64), .Y(ab_18__4_) );
  AND2X1_RVT U475 ( .A1(n27), .A2(n61), .Y(ab_18__3_) );
  AND2X1_RVT U476 ( .A1(n27), .A2(n59), .Y(ab_18__2_) );
  AND2X1_RVT U477 ( .A1(A[18]), .A2(n57), .Y(ab_18__1_) );
  AND2X1_RVT U478 ( .A1(n27), .A2(n8), .Y(ab_18__13_) );
  AND2X1_RVT U479 ( .A1(n27), .A2(n7), .Y(ab_18__12_) );
  AND2X1_RVT U480 ( .A1(n27), .A2(n6), .Y(ab_18__11_) );
  AND2X1_RVT U481 ( .A1(n27), .A2(n3), .Y(ab_18__10_) );
  AND2X1_RVT U482 ( .A1(n27), .A2(n56), .Y(ab_18__0_) );
  AND2X1_RVT U483 ( .A1(n26), .A2(n74), .Y(ab_17__9_) );
  AND2X1_RVT U484 ( .A1(n26), .A2(n72), .Y(ab_17__8_) );
  AND2X1_RVT U485 ( .A1(n26), .A2(n70), .Y(ab_17__7_) );
  AND2X1_RVT U486 ( .A1(n26), .A2(n68), .Y(ab_17__6_) );
  AND2X1_RVT U487 ( .A1(n26), .A2(n66), .Y(ab_17__5_) );
  AND2X1_RVT U488 ( .A1(n26), .A2(n64), .Y(ab_17__4_) );
  AND2X1_RVT U489 ( .A1(n26), .A2(n61), .Y(ab_17__3_) );
  AND2X1_RVT U490 ( .A1(n26), .A2(n59), .Y(ab_17__2_) );
  AND2X1_RVT U491 ( .A1(A[17]), .A2(n57), .Y(ab_17__1_) );
  AND2X1_RVT U492 ( .A1(n26), .A2(B[14]), .Y(ab_17__14_) );
  AND2X1_RVT U493 ( .A1(n26), .A2(n8), .Y(ab_17__13_) );
  AND2X1_RVT U494 ( .A1(n26), .A2(B[12]), .Y(ab_17__12_) );
  AND2X1_RVT U495 ( .A1(n26), .A2(n6), .Y(ab_17__11_) );
  AND2X1_RVT U496 ( .A1(n26), .A2(n4), .Y(ab_17__10_) );
  AND2X1_RVT U497 ( .A1(A[17]), .A2(n56), .Y(ab_17__0_) );
  AND2X1_RVT U498 ( .A1(n25), .A2(n74), .Y(ab_16__9_) );
  AND2X1_RVT U499 ( .A1(n25), .A2(n72), .Y(ab_16__8_) );
  AND2X1_RVT U500 ( .A1(n25), .A2(n70), .Y(ab_16__7_) );
  AND2X1_RVT U501 ( .A1(n25), .A2(n68), .Y(ab_16__6_) );
  AND2X1_RVT U502 ( .A1(n25), .A2(n66), .Y(ab_16__5_) );
  AND2X1_RVT U503 ( .A1(n25), .A2(n64), .Y(ab_16__4_) );
  AND2X1_RVT U504 ( .A1(A[16]), .A2(n61), .Y(ab_16__3_) );
  AND2X1_RVT U505 ( .A1(n25), .A2(n59), .Y(ab_16__2_) );
  AND2X1_RVT U506 ( .A1(A[16]), .A2(n57), .Y(ab_16__1_) );
  AND2X1_RVT U507 ( .A1(n25), .A2(n10), .Y(ab_16__15_) );
  AND2X1_RVT U508 ( .A1(n25), .A2(n9), .Y(ab_16__14_) );
  AND2X1_RVT U509 ( .A1(n25), .A2(n8), .Y(ab_16__13_) );
  AND2X1_RVT U510 ( .A1(n25), .A2(n7), .Y(ab_16__12_) );
  AND2X1_RVT U511 ( .A1(n25), .A2(n6), .Y(ab_16__11_) );
  AND2X1_RVT U512 ( .A1(n25), .A2(n3), .Y(ab_16__10_) );
  AND2X1_RVT U513 ( .A1(n25), .A2(n56), .Y(ab_16__0_) );
  AND2X1_RVT U514 ( .A1(n24), .A2(n74), .Y(ab_15__9_) );
  AND2X1_RVT U515 ( .A1(n24), .A2(n72), .Y(ab_15__8_) );
  AND2X1_RVT U516 ( .A1(n24), .A2(n70), .Y(ab_15__7_) );
  AND2X1_RVT U517 ( .A1(n24), .A2(n68), .Y(ab_15__6_) );
  AND2X1_RVT U518 ( .A1(n24), .A2(n66), .Y(ab_15__5_) );
  AND2X1_RVT U519 ( .A1(n24), .A2(n64), .Y(ab_15__4_) );
  AND2X1_RVT U520 ( .A1(A[15]), .A2(n61), .Y(ab_15__3_) );
  AND2X1_RVT U521 ( .A1(n24), .A2(n59), .Y(ab_15__2_) );
  AND2X1_RVT U522 ( .A1(A[15]), .A2(n57), .Y(ab_15__1_) );
  AND2X1_RVT U523 ( .A1(n24), .A2(n11), .Y(ab_15__16_) );
  AND2X1_RVT U524 ( .A1(n24), .A2(n10), .Y(ab_15__15_) );
  AND2X1_RVT U525 ( .A1(n24), .A2(B[14]), .Y(ab_15__14_) );
  AND2X1_RVT U526 ( .A1(n24), .A2(n8), .Y(ab_15__13_) );
  AND2X1_RVT U527 ( .A1(n24), .A2(B[12]), .Y(ab_15__12_) );
  AND2X1_RVT U528 ( .A1(n24), .A2(n6), .Y(ab_15__11_) );
  AND2X1_RVT U529 ( .A1(n24), .A2(n4), .Y(ab_15__10_) );
  AND2X1_RVT U530 ( .A1(A[15]), .A2(n56), .Y(ab_15__0_) );
  AND2X1_RVT U531 ( .A1(n23), .A2(n74), .Y(ab_14__9_) );
  AND2X1_RVT U532 ( .A1(n23), .A2(n72), .Y(ab_14__8_) );
  AND2X1_RVT U533 ( .A1(n23), .A2(n70), .Y(ab_14__7_) );
  AND2X1_RVT U534 ( .A1(n23), .A2(n68), .Y(ab_14__6_) );
  AND2X1_RVT U535 ( .A1(n23), .A2(n66), .Y(ab_14__5_) );
  AND2X1_RVT U536 ( .A1(A[14]), .A2(n64), .Y(ab_14__4_) );
  AND2X1_RVT U537 ( .A1(n23), .A2(n61), .Y(ab_14__3_) );
  AND2X1_RVT U538 ( .A1(A[14]), .A2(n59), .Y(ab_14__2_) );
  AND2X1_RVT U539 ( .A1(n23), .A2(n57), .Y(ab_14__1_) );
  AND2X1_RVT U540 ( .A1(A[14]), .A2(n12), .Y(ab_14__17_) );
  AND2X1_RVT U541 ( .A1(n23), .A2(B[16]), .Y(ab_14__16_) );
  AND2X1_RVT U542 ( .A1(n23), .A2(n10), .Y(ab_14__15_) );
  AND2X1_RVT U543 ( .A1(n23), .A2(n9), .Y(ab_14__14_) );
  AND2X1_RVT U544 ( .A1(n23), .A2(n8), .Y(ab_14__13_) );
  AND2X1_RVT U545 ( .A1(n23), .A2(n7), .Y(ab_14__12_) );
  AND2X1_RVT U546 ( .A1(n23), .A2(n6), .Y(ab_14__11_) );
  AND2X1_RVT U547 ( .A1(n23), .A2(n3), .Y(ab_14__10_) );
  AND2X1_RVT U548 ( .A1(A[14]), .A2(n56), .Y(ab_14__0_) );
  AND2X1_RVT U549 ( .A1(n22), .A2(n74), .Y(ab_13__9_) );
  AND2X1_RVT U550 ( .A1(n22), .A2(n72), .Y(ab_13__8_) );
  AND2X1_RVT U551 ( .A1(A[13]), .A2(n70), .Y(ab_13__7_) );
  AND2X1_RVT U552 ( .A1(n22), .A2(n68), .Y(ab_13__6_) );
  AND2X1_RVT U553 ( .A1(A[13]), .A2(n66), .Y(ab_13__5_) );
  AND2X1_RVT U554 ( .A1(n22), .A2(n64), .Y(ab_13__4_) );
  AND2X1_RVT U555 ( .A1(A[13]), .A2(n61), .Y(ab_13__3_) );
  AND2X1_RVT U556 ( .A1(n22), .A2(n59), .Y(ab_13__2_) );
  AND2X1_RVT U557 ( .A1(A[13]), .A2(n57), .Y(ab_13__1_) );
  AND2X1_RVT U558 ( .A1(n22), .A2(n13), .Y(ab_13__18_) );
  AND2X1_RVT U559 ( .A1(n22), .A2(n12), .Y(ab_13__17_) );
  AND2X1_RVT U560 ( .A1(n22), .A2(n11), .Y(ab_13__16_) );
  AND2X1_RVT U561 ( .A1(n22), .A2(n10), .Y(ab_13__15_) );
  AND2X1_RVT U562 ( .A1(n22), .A2(B[14]), .Y(ab_13__14_) );
  AND2X1_RVT U563 ( .A1(n22), .A2(n8), .Y(ab_13__13_) );
  AND2X1_RVT U564 ( .A1(n22), .A2(B[12]), .Y(ab_13__12_) );
  AND2X1_RVT U565 ( .A1(n22), .A2(n6), .Y(ab_13__11_) );
  AND2X1_RVT U566 ( .A1(n22), .A2(n4), .Y(ab_13__10_) );
  AND2X1_RVT U567 ( .A1(A[13]), .A2(n56), .Y(ab_13__0_) );
  AND2X1_RVT U568 ( .A1(n21), .A2(n74), .Y(ab_12__9_) );
  AND2X1_RVT U569 ( .A1(n21), .A2(n72), .Y(ab_12__8_) );
  AND2X1_RVT U570 ( .A1(n21), .A2(n70), .Y(ab_12__7_) );
  AND2X1_RVT U571 ( .A1(A[12]), .A2(n68), .Y(ab_12__6_) );
  AND2X1_RVT U572 ( .A1(n21), .A2(n66), .Y(ab_12__5_) );
  AND2X1_RVT U573 ( .A1(A[12]), .A2(n64), .Y(ab_12__4_) );
  AND2X1_RVT U574 ( .A1(n21), .A2(n61), .Y(ab_12__3_) );
  AND2X1_RVT U575 ( .A1(A[12]), .A2(n59), .Y(ab_12__2_) );
  AND2X1_RVT U576 ( .A1(n21), .A2(n58), .Y(ab_12__1_) );
  AND2X1_RVT U577 ( .A1(A[12]), .A2(n15), .Y(ab_12__19_) );
  AND2X1_RVT U578 ( .A1(n21), .A2(n13), .Y(ab_12__18_) );
  AND2X1_RVT U579 ( .A1(n21), .A2(n12), .Y(ab_12__17_) );
  AND2X1_RVT U580 ( .A1(n21), .A2(n11), .Y(ab_12__16_) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n10), .Y(ab_12__15_) );
  AND2X1_RVT U582 ( .A1(n21), .A2(n9), .Y(ab_12__14_) );
  AND2X1_RVT U583 ( .A1(n21), .A2(n8), .Y(ab_12__13_) );
  AND2X1_RVT U584 ( .A1(n21), .A2(n7), .Y(ab_12__12_) );
  AND2X1_RVT U585 ( .A1(n21), .A2(n6), .Y(ab_12__11_) );
  AND2X1_RVT U586 ( .A1(n21), .A2(n3), .Y(ab_12__10_) );
  AND2X1_RVT U587 ( .A1(A[12]), .A2(n56), .Y(ab_12__0_) );
  AND2X1_RVT U588 ( .A1(n20), .A2(n74), .Y(ab_11__9_) );
  AND2X1_RVT U589 ( .A1(n20), .A2(n72), .Y(ab_11__8_) );
  AND2X1_RVT U590 ( .A1(A[11]), .A2(n70), .Y(ab_11__7_) );
  AND2X1_RVT U591 ( .A1(n20), .A2(n68), .Y(ab_11__6_) );
  AND2X1_RVT U592 ( .A1(A[11]), .A2(n66), .Y(ab_11__5_) );
  AND2X1_RVT U593 ( .A1(n20), .A2(n64), .Y(ab_11__4_) );
  AND2X1_RVT U594 ( .A1(A[11]), .A2(n61), .Y(ab_11__3_) );
  AND2X1_RVT U595 ( .A1(n20), .A2(n60), .Y(ab_11__2_) );
  AND2X1_RVT U596 ( .A1(A[11]), .A2(n17), .Y(ab_11__20_) );
  AND2X1_RVT U597 ( .A1(n20), .A2(n58), .Y(ab_11__1_) );
  AND2X1_RVT U598 ( .A1(A[11]), .A2(n15), .Y(ab_11__19_) );
  AND2X1_RVT U599 ( .A1(n20), .A2(n13), .Y(ab_11__18_) );
  AND2X1_RVT U600 ( .A1(n20), .A2(n12), .Y(ab_11__17_) );
  AND2X1_RVT U601 ( .A1(n20), .A2(n11), .Y(ab_11__16_) );
  AND2X1_RVT U602 ( .A1(n20), .A2(n10), .Y(ab_11__15_) );
  AND2X1_RVT U603 ( .A1(n20), .A2(n9), .Y(ab_11__14_) );
  AND2X1_RVT U604 ( .A1(n20), .A2(n8), .Y(ab_11__13_) );
  AND2X1_RVT U605 ( .A1(n20), .A2(n7), .Y(ab_11__12_) );
  AND2X1_RVT U606 ( .A1(n20), .A2(n6), .Y(ab_11__11_) );
  AND2X1_RVT U607 ( .A1(n20), .A2(n4), .Y(ab_11__10_) );
  AND2X1_RVT U608 ( .A1(A[11]), .A2(n56), .Y(ab_11__0_) );
  AND2X1_RVT U609 ( .A1(n18), .A2(n74), .Y(ab_10__9_) );
  AND2X1_RVT U610 ( .A1(n19), .A2(n72), .Y(ab_10__8_) );
  AND2X1_RVT U611 ( .A1(n18), .A2(n70), .Y(ab_10__7_) );
  AND2X1_RVT U612 ( .A1(n19), .A2(n68), .Y(ab_10__6_) );
  AND2X1_RVT U613 ( .A1(n18), .A2(n66), .Y(ab_10__5_) );
  AND2X1_RVT U614 ( .A1(n19), .A2(n64), .Y(ab_10__4_) );
  AND2X1_RVT U615 ( .A1(n18), .A2(n62), .Y(ab_10__3_) );
  AND2X1_RVT U616 ( .A1(n19), .A2(n60), .Y(ab_10__2_) );
  AND2X1_RVT U617 ( .A1(n18), .A2(B[21]), .Y(ab_10__21_) );
  AND2X1_RVT U618 ( .A1(n19), .A2(n17), .Y(ab_10__20_) );
  AND2X1_RVT U619 ( .A1(n18), .A2(n58), .Y(ab_10__1_) );
  AND2X1_RVT U620 ( .A1(n19), .A2(n15), .Y(ab_10__19_) );
  AND2X1_RVT U621 ( .A1(n18), .A2(n13), .Y(ab_10__18_) );
  AND2X1_RVT U622 ( .A1(n19), .A2(n12), .Y(ab_10__17_) );
  AND2X1_RVT U623 ( .A1(n18), .A2(n11), .Y(ab_10__16_) );
  AND2X1_RVT U624 ( .A1(n19), .A2(n10), .Y(ab_10__15_) );
  AND2X1_RVT U625 ( .A1(n18), .A2(n9), .Y(ab_10__14_) );
  AND2X1_RVT U626 ( .A1(n19), .A2(n8), .Y(ab_10__13_) );
  AND2X1_RVT U627 ( .A1(n18), .A2(n7), .Y(ab_10__12_) );
  AND2X1_RVT U628 ( .A1(n19), .A2(n6), .Y(ab_10__11_) );
  AND2X1_RVT U629 ( .A1(n18), .A2(n3), .Y(ab_10__10_) );
  AND2X1_RVT U630 ( .A1(n19), .A2(n56), .Y(ab_10__0_) );
  AND2X1_RVT U631 ( .A1(n35), .A2(n74), .Y(ab_0__9_) );
  AND2X1_RVT U632 ( .A1(n35), .A2(n72), .Y(ab_0__8_) );
  AND2X1_RVT U633 ( .A1(n35), .A2(n70), .Y(ab_0__7_) );
  AND2X1_RVT U634 ( .A1(n35), .A2(n68), .Y(ab_0__6_) );
  AND2X1_RVT U635 ( .A1(n35), .A2(n66), .Y(ab_0__5_) );
  AND2X1_RVT U636 ( .A1(n35), .A2(n63), .Y(ab_0__4_) );
  AND2X1_RVT U637 ( .A1(n35), .A2(n62), .Y(ab_0__3_) );
  AND2X1_RVT U638 ( .A1(n35), .A2(B[31]), .Y(ab_0__31_) );
  AND2X1_RVT U639 ( .A1(n34), .A2(B[30]), .Y(ab_0__30_) );
  AND2X1_RVT U640 ( .A1(n34), .A2(n60), .Y(ab_0__2_) );
  AND2X1_RVT U641 ( .A1(n34), .A2(B[29]), .Y(ab_0__29_) );
  AND2X1_RVT U642 ( .A1(n34), .A2(B[28]), .Y(ab_0__28_) );
  AND2X1_RVT U643 ( .A1(n34), .A2(B[27]), .Y(ab_0__27_) );
  AND2X1_RVT U644 ( .A1(n34), .A2(B[26]), .Y(ab_0__26_) );
  AND2X1_RVT U645 ( .A1(n34), .A2(B[25]), .Y(ab_0__25_) );
  AND2X1_RVT U646 ( .A1(n34), .A2(B[24]), .Y(ab_0__24_) );
  AND2X1_RVT U647 ( .A1(n34), .A2(B[23]), .Y(ab_0__23_) );
  AND2X1_RVT U648 ( .A1(n34), .A2(B[22]), .Y(ab_0__22_) );
  AND2X1_RVT U649 ( .A1(n34), .A2(B[21]), .Y(ab_0__21_) );
  AND2X1_RVT U650 ( .A1(n34), .A2(B[20]), .Y(ab_0__20_) );
  AND2X1_RVT U651 ( .A1(n33), .A2(n58), .Y(ab_0__1_) );
  AND2X1_RVT U652 ( .A1(n33), .A2(B[19]), .Y(ab_0__19_) );
  AND2X1_RVT U653 ( .A1(n33), .A2(n13), .Y(ab_0__18_) );
  AND2X1_RVT U654 ( .A1(n33), .A2(n12), .Y(ab_0__17_) );
  AND2X1_RVT U655 ( .A1(n33), .A2(n11), .Y(ab_0__16_) );
  AND2X1_RVT U656 ( .A1(n33), .A2(B[15]), .Y(ab_0__15_) );
  AND2X1_RVT U657 ( .A1(n33), .A2(n9), .Y(ab_0__14_) );
  AND2X1_RVT U658 ( .A1(n33), .A2(n8), .Y(ab_0__13_) );
  AND2X1_RVT U659 ( .A1(n33), .A2(n7), .Y(ab_0__12_) );
  AND2X1_RVT U660 ( .A1(n33), .A2(n6), .Y(ab_0__11_) );
  AND2X1_RVT U661 ( .A1(n33), .A2(n4), .Y(ab_0__10_) );
  AND2X1_RVT U662 ( .A1(n33), .A2(n56), .Y(PRODUCT_0_) );
endmodule


module OSPE_1_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;

  wire   [31:1] carry;

  FADDX1_RVT U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1_RVT U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1_RVT U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1_RVT U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1_RVT U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1_RVT U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1_RVT U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1_RVT U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module OSPE_1 ( clk, rstnPipe, rstnPsum, ipA, ipB, opA, opB, opC );
  input [31:0] ipA;
  input [31:0] ipB;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] opC;
  input clk, rstnPipe, rstnPsum;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N9, N8, N7, N6, N5, N4, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n1, n2, n3, n4, n5, n6,
         n7;
  wire   [31:0] opC_wire;

  AND2X1_RVT U3 ( .A1(n1), .A2(ipB[30]), .Y(N99) );
  AND2X1_RVT U4 ( .A1(ipB[29]), .A2(n1), .Y(N98) );
  AND2X1_RVT U5 ( .A1(ipB[28]), .A2(n1), .Y(N97) );
  AND2X1_RVT U6 ( .A1(ipB[27]), .A2(n1), .Y(N96) );
  AND2X1_RVT U7 ( .A1(ipB[26]), .A2(n1), .Y(N95) );
  AND2X1_RVT U8 ( .A1(ipB[25]), .A2(n1), .Y(N94) );
  AND2X1_RVT U9 ( .A1(ipB[24]), .A2(n1), .Y(N93) );
  AND2X1_RVT U10 ( .A1(ipB[23]), .A2(n1), .Y(N92) );
  AND2X1_RVT U11 ( .A1(ipB[22]), .A2(n1), .Y(N91) );
  AND2X1_RVT U12 ( .A1(ipB[21]), .A2(n1), .Y(N90) );
  AND2X1_RVT U13 ( .A1(ipB[20]), .A2(n1), .Y(N89) );
  AND2X1_RVT U14 ( .A1(ipB[19]), .A2(n1), .Y(N88) );
  AND2X1_RVT U15 ( .A1(ipB[18]), .A2(n1), .Y(N87) );
  AND2X1_RVT U16 ( .A1(ipB[17]), .A2(n2), .Y(N86) );
  AND2X1_RVT U17 ( .A1(ipB[16]), .A2(n2), .Y(N85) );
  AND2X1_RVT U18 ( .A1(ipB[15]), .A2(n2), .Y(N84) );
  AND2X1_RVT U19 ( .A1(ipB[14]), .A2(n2), .Y(N83) );
  AND2X1_RVT U20 ( .A1(ipB[13]), .A2(n2), .Y(N82) );
  AND2X1_RVT U21 ( .A1(ipB[12]), .A2(n2), .Y(N81) );
  AND2X1_RVT U22 ( .A1(ipB[11]), .A2(n2), .Y(N80) );
  AND2X1_RVT U23 ( .A1(ipB[10]), .A2(n2), .Y(N79) );
  AND2X1_RVT U24 ( .A1(ipB[9]), .A2(n2), .Y(N78) );
  AND2X1_RVT U25 ( .A1(ipB[8]), .A2(n2), .Y(N77) );
  AND2X1_RVT U26 ( .A1(ipB[7]), .A2(n2), .Y(N76) );
  AND2X1_RVT U27 ( .A1(ipB[6]), .A2(n2), .Y(N75) );
  AND2X1_RVT U28 ( .A1(ipB[5]), .A2(n2), .Y(N74) );
  AND2X1_RVT U29 ( .A1(ipB[4]), .A2(n2), .Y(N73) );
  AND2X1_RVT U30 ( .A1(ipB[3]), .A2(n3), .Y(N72) );
  AND2X1_RVT U31 ( .A1(ipB[2]), .A2(n3), .Y(N71) );
  AND2X1_RVT U32 ( .A1(ipB[1]), .A2(n3), .Y(N70) );
  AND2X1_RVT U33 ( .A1(ipB[0]), .A2(n3), .Y(N69) );
  AND2X1_RVT U34 ( .A1(ipA[31]), .A2(n3), .Y(N68) );
  AND2X1_RVT U35 ( .A1(ipA[30]), .A2(n3), .Y(N67) );
  AND2X1_RVT U36 ( .A1(ipA[29]), .A2(n3), .Y(N66) );
  AND2X1_RVT U37 ( .A1(ipA[28]), .A2(n3), .Y(N65) );
  AND2X1_RVT U38 ( .A1(ipA[27]), .A2(n3), .Y(N64) );
  AND2X1_RVT U39 ( .A1(ipA[26]), .A2(n3), .Y(N63) );
  AND2X1_RVT U40 ( .A1(ipA[25]), .A2(n3), .Y(N62) );
  AND2X1_RVT U41 ( .A1(ipA[24]), .A2(n3), .Y(N61) );
  AND2X1_RVT U42 ( .A1(ipA[23]), .A2(n3), .Y(N60) );
  AND2X1_RVT U43 ( .A1(ipA[22]), .A2(n3), .Y(N59) );
  AND2X1_RVT U44 ( .A1(ipA[21]), .A2(n4), .Y(N58) );
  AND2X1_RVT U45 ( .A1(ipA[20]), .A2(n4), .Y(N57) );
  AND2X1_RVT U46 ( .A1(ipA[19]), .A2(n4), .Y(N56) );
  AND2X1_RVT U47 ( .A1(ipA[18]), .A2(n4), .Y(N55) );
  AND2X1_RVT U48 ( .A1(ipA[17]), .A2(n4), .Y(N54) );
  AND2X1_RVT U49 ( .A1(ipA[16]), .A2(n4), .Y(N53) );
  AND2X1_RVT U50 ( .A1(ipA[15]), .A2(n4), .Y(N52) );
  AND2X1_RVT U51 ( .A1(ipA[14]), .A2(n4), .Y(N51) );
  AND2X1_RVT U52 ( .A1(ipA[13]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(ipA[12]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(ipA[11]), .A2(n4), .Y(N48) );
  AND2X1_RVT U55 ( .A1(ipA[10]), .A2(n4), .Y(N47) );
  AND2X1_RVT U56 ( .A1(ipA[9]), .A2(n4), .Y(N46) );
  AND2X1_RVT U57 ( .A1(ipA[8]), .A2(n4), .Y(N45) );
  AND2X1_RVT U58 ( .A1(ipA[7]), .A2(n5), .Y(N44) );
  AND2X1_RVT U59 ( .A1(ipA[6]), .A2(n5), .Y(N43) );
  AND2X1_RVT U60 ( .A1(ipA[5]), .A2(n5), .Y(N42) );
  AND2X1_RVT U61 ( .A1(ipA[4]), .A2(n5), .Y(N41) );
  AND2X1_RVT U62 ( .A1(ipA[3]), .A2(n5), .Y(N40) );
  AND2X1_RVT U63 ( .A1(ipA[2]), .A2(n5), .Y(N39) );
  AND2X1_RVT U64 ( .A1(ipA[1]), .A2(n5), .Y(N38) );
  AND2X1_RVT U65 ( .A1(ipA[0]), .A2(n5), .Y(N37) );
  AND2X1_RVT U66 ( .A1(n6), .A2(opC_wire[31]), .Y(N133) );
  AND2X1_RVT U67 ( .A1(opC_wire[30]), .A2(n7), .Y(N132) );
  AND2X1_RVT U68 ( .A1(opC_wire[29]), .A2(n6), .Y(N131) );
  AND2X1_RVT U69 ( .A1(opC_wire[28]), .A2(n7), .Y(N130) );
  AND2X1_RVT U70 ( .A1(opC_wire[27]), .A2(n7), .Y(N129) );
  AND2X1_RVT U71 ( .A1(opC_wire[26]), .A2(n7), .Y(N128) );
  AND2X1_RVT U72 ( .A1(opC_wire[25]), .A2(n7), .Y(N127) );
  AND2X1_RVT U73 ( .A1(opC_wire[24]), .A2(n7), .Y(N126) );
  AND2X1_RVT U74 ( .A1(opC_wire[23]), .A2(n7), .Y(N125) );
  AND2X1_RVT U75 ( .A1(opC_wire[22]), .A2(n7), .Y(N124) );
  AND2X1_RVT U76 ( .A1(opC_wire[21]), .A2(n7), .Y(N123) );
  AND2X1_RVT U77 ( .A1(opC_wire[20]), .A2(n7), .Y(N122) );
  AND2X1_RVT U78 ( .A1(opC_wire[19]), .A2(n7), .Y(N121) );
  AND2X1_RVT U79 ( .A1(opC_wire[18]), .A2(n6), .Y(N120) );
  AND2X1_RVT U80 ( .A1(opC_wire[17]), .A2(n6), .Y(N119) );
  AND2X1_RVT U81 ( .A1(opC_wire[16]), .A2(n6), .Y(N118) );
  AND2X1_RVT U82 ( .A1(opC_wire[15]), .A2(n6), .Y(N117) );
  AND2X1_RVT U83 ( .A1(opC_wire[14]), .A2(n6), .Y(N116) );
  AND2X1_RVT U84 ( .A1(opC_wire[13]), .A2(n6), .Y(N115) );
  AND2X1_RVT U85 ( .A1(opC_wire[12]), .A2(n6), .Y(N114) );
  AND2X1_RVT U86 ( .A1(opC_wire[11]), .A2(n6), .Y(N113) );
  AND2X1_RVT U87 ( .A1(opC_wire[10]), .A2(n6), .Y(N112) );
  AND2X1_RVT U88 ( .A1(opC_wire[9]), .A2(n6), .Y(N111) );
  AND2X1_RVT U89 ( .A1(opC_wire[8]), .A2(n6), .Y(N110) );
  AND2X1_RVT U90 ( .A1(opC_wire[7]), .A2(n6), .Y(N109) );
  AND2X1_RVT U91 ( .A1(opC_wire[6]), .A2(n6), .Y(N108) );
  AND2X1_RVT U92 ( .A1(opC_wire[5]), .A2(n6), .Y(N107) );
  AND2X1_RVT U93 ( .A1(opC_wire[4]), .A2(n7), .Y(N106) );
  AND2X1_RVT U94 ( .A1(opC_wire[3]), .A2(n7), .Y(N105) );
  AND2X1_RVT U95 ( .A1(opC_wire[2]), .A2(n7), .Y(N104) );
  AND2X1_RVT U96 ( .A1(opC_wire[1]), .A2(n7), .Y(N103) );
  AND2X1_RVT U97 ( .A1(opC_wire[0]), .A2(n7), .Y(N102) );
  AND2X1_RVT U98 ( .A1(ipB[31]), .A2(n5), .Y(N100) );
  OSPE_1_DW02_mult_0 mult_23 ( .A(ipA), .B(ipB), .PRODUCT_31_(N35), 
        .PRODUCT_30_(N34), .PRODUCT_29_(N33), .PRODUCT_28_(N32), .PRODUCT_27_(
        N31), .PRODUCT_26_(N30), .PRODUCT_25_(N29), .PRODUCT_24_(N28), 
        .PRODUCT_23_(N27), .PRODUCT_22_(N26), .PRODUCT_21_(N25), .PRODUCT_20_(
        N24), .PRODUCT_19_(N23), .PRODUCT_18_(N22), .PRODUCT_17_(N21), 
        .PRODUCT_16_(N20), .PRODUCT_15_(N19), .PRODUCT_14_(N18), .PRODUCT_13_(
        N17), .PRODUCT_12_(N16), .PRODUCT_11_(N15), .PRODUCT_10_(N14), 
        .PRODUCT_9_(N13), .PRODUCT_8_(N12), .PRODUCT_7_(N11), .PRODUCT_6_(N10), 
        .PRODUCT_5_(N9), .PRODUCT_4_(N8), .PRODUCT_3_(N7), .PRODUCT_2_(N6), 
        .PRODUCT_1_(N5), .PRODUCT_0_(N4) );
  OSPE_1_DW01_add_0 add_23 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4}), .B(opC), .SUM(opC_wire) );
  DFFX1_RVT opC_reg_31_ ( .D(N133), .CLK(clk), .Q(opC[31]) );
  DFFX1_RVT opC_reg_30_ ( .D(N132), .CLK(clk), .Q(opC[30]) );
  DFFX1_RVT opC_reg_29_ ( .D(N131), .CLK(clk), .Q(opC[29]) );
  DFFX1_RVT opC_reg_28_ ( .D(N130), .CLK(clk), .Q(opC[28]) );
  DFFX1_RVT opC_reg_27_ ( .D(N129), .CLK(clk), .Q(opC[27]) );
  DFFX1_RVT opC_reg_26_ ( .D(N128), .CLK(clk), .Q(opC[26]) );
  DFFX1_RVT opC_reg_25_ ( .D(N127), .CLK(clk), .Q(opC[25]) );
  DFFX1_RVT opC_reg_24_ ( .D(N126), .CLK(clk), .Q(opC[24]) );
  DFFX1_RVT opC_reg_23_ ( .D(N125), .CLK(clk), .Q(opC[23]) );
  DFFX1_RVT opC_reg_22_ ( .D(N124), .CLK(clk), .Q(opC[22]) );
  DFFX1_RVT opC_reg_21_ ( .D(N123), .CLK(clk), .Q(opC[21]) );
  DFFX1_RVT opC_reg_20_ ( .D(N122), .CLK(clk), .Q(opC[20]) );
  DFFX1_RVT opC_reg_19_ ( .D(N121), .CLK(clk), .Q(opC[19]) );
  DFFX1_RVT opC_reg_18_ ( .D(N120), .CLK(clk), .Q(opC[18]) );
  DFFX1_RVT opC_reg_17_ ( .D(N119), .CLK(clk), .Q(opC[17]) );
  DFFX1_RVT opC_reg_16_ ( .D(N118), .CLK(clk), .Q(opC[16]) );
  DFFX1_RVT opC_reg_15_ ( .D(N117), .CLK(clk), .Q(opC[15]) );
  DFFX1_RVT opC_reg_14_ ( .D(N116), .CLK(clk), .Q(opC[14]) );
  DFFX1_RVT opC_reg_13_ ( .D(N115), .CLK(clk), .Q(opC[13]) );
  DFFX1_RVT opC_reg_12_ ( .D(N114), .CLK(clk), .Q(opC[12]) );
  DFFX1_RVT opC_reg_11_ ( .D(N113), .CLK(clk), .Q(opC[11]) );
  DFFX1_RVT opC_reg_10_ ( .D(N112), .CLK(clk), .Q(opC[10]) );
  DFFX1_RVT opC_reg_9_ ( .D(N111), .CLK(clk), .Q(opC[9]) );
  DFFX1_RVT opC_reg_8_ ( .D(N110), .CLK(clk), .Q(opC[8]) );
  DFFX1_RVT opC_reg_7_ ( .D(N109), .CLK(clk), .Q(opC[7]) );
  DFFX1_RVT opC_reg_6_ ( .D(N108), .CLK(clk), .Q(opC[6]) );
  DFFX1_RVT opC_reg_0_ ( .D(N102), .CLK(clk), .Q(opC[0]) );
  DFFX1_RVT opC_reg_5_ ( .D(N107), .CLK(clk), .Q(opC[5]) );
  DFFX1_RVT opC_reg_4_ ( .D(N106), .CLK(clk), .Q(opC[4]) );
  DFFX1_RVT opC_reg_3_ ( .D(N105), .CLK(clk), .Q(opC[3]) );
  DFFX1_RVT opC_reg_2_ ( .D(N104), .CLK(clk), .Q(opC[2]) );
  DFFX1_RVT opC_reg_1_ ( .D(N103), .CLK(clk), .Q(opC[1]) );
  DFFX1_RVT opA_reg_31_ ( .D(N68), .CLK(clk), .Q(opA[31]) );
  DFFX1_RVT opA_reg_30_ ( .D(N67), .CLK(clk), .Q(opA[30]) );
  DFFX1_RVT opA_reg_29_ ( .D(N66), .CLK(clk), .Q(opA[29]) );
  DFFX1_RVT opA_reg_28_ ( .D(N65), .CLK(clk), .Q(opA[28]) );
  DFFX1_RVT opA_reg_27_ ( .D(N64), .CLK(clk), .Q(opA[27]) );
  DFFX1_RVT opA_reg_26_ ( .D(N63), .CLK(clk), .Q(opA[26]) );
  DFFX1_RVT opA_reg_25_ ( .D(N62), .CLK(clk), .Q(opA[25]) );
  DFFX1_RVT opA_reg_24_ ( .D(N61), .CLK(clk), .Q(opA[24]) );
  DFFX1_RVT opA_reg_23_ ( .D(N60), .CLK(clk), .Q(opA[23]) );
  DFFX1_RVT opA_reg_22_ ( .D(N59), .CLK(clk), .Q(opA[22]) );
  DFFX1_RVT opA_reg_21_ ( .D(N58), .CLK(clk), .Q(opA[21]) );
  DFFX1_RVT opA_reg_20_ ( .D(N57), .CLK(clk), .Q(opA[20]) );
  DFFX1_RVT opA_reg_19_ ( .D(N56), .CLK(clk), .Q(opA[19]) );
  DFFX1_RVT opA_reg_18_ ( .D(N55), .CLK(clk), .Q(opA[18]) );
  DFFX1_RVT opA_reg_17_ ( .D(N54), .CLK(clk), .Q(opA[17]) );
  DFFX1_RVT opA_reg_16_ ( .D(N53), .CLK(clk), .Q(opA[16]) );
  DFFX1_RVT opA_reg_15_ ( .D(N52), .CLK(clk), .Q(opA[15]) );
  DFFX1_RVT opA_reg_14_ ( .D(N51), .CLK(clk), .Q(opA[14]) );
  DFFX1_RVT opA_reg_13_ ( .D(N50), .CLK(clk), .Q(opA[13]) );
  DFFX1_RVT opA_reg_12_ ( .D(N49), .CLK(clk), .Q(opA[12]) );
  DFFX1_RVT opA_reg_11_ ( .D(N48), .CLK(clk), .Q(opA[11]) );
  DFFX1_RVT opA_reg_10_ ( .D(N47), .CLK(clk), .Q(opA[10]) );
  DFFX1_RVT opA_reg_9_ ( .D(N46), .CLK(clk), .Q(opA[9]) );
  DFFX1_RVT opA_reg_8_ ( .D(N45), .CLK(clk), .Q(opA[8]) );
  DFFX1_RVT opA_reg_7_ ( .D(N44), .CLK(clk), .Q(opA[7]) );
  DFFX1_RVT opA_reg_6_ ( .D(N43), .CLK(clk), .Q(opA[6]) );
  DFFX1_RVT opA_reg_5_ ( .D(N42), .CLK(clk), .Q(opA[5]) );
  DFFX1_RVT opA_reg_4_ ( .D(N41), .CLK(clk), .Q(opA[4]) );
  DFFX1_RVT opA_reg_3_ ( .D(N40), .CLK(clk), .Q(opA[3]) );
  DFFX1_RVT opA_reg_2_ ( .D(N39), .CLK(clk), .Q(opA[2]) );
  DFFX1_RVT opA_reg_1_ ( .D(N38), .CLK(clk), .Q(opA[1]) );
  DFFX1_RVT opA_reg_0_ ( .D(N37), .CLK(clk), .Q(opA[0]) );
  DFFX1_RVT opB_reg_31_ ( .D(N100), .CLK(clk), .Q(opB[31]) );
  DFFX1_RVT opB_reg_30_ ( .D(N99), .CLK(clk), .Q(opB[30]) );
  DFFX1_RVT opB_reg_29_ ( .D(N98), .CLK(clk), .Q(opB[29]) );
  DFFX1_RVT opB_reg_28_ ( .D(N97), .CLK(clk), .Q(opB[28]) );
  DFFX1_RVT opB_reg_27_ ( .D(N96), .CLK(clk), .Q(opB[27]) );
  DFFX1_RVT opB_reg_26_ ( .D(N95), .CLK(clk), .Q(opB[26]) );
  DFFX1_RVT opB_reg_25_ ( .D(N94), .CLK(clk), .Q(opB[25]) );
  DFFX1_RVT opB_reg_24_ ( .D(N93), .CLK(clk), .Q(opB[24]) );
  DFFX1_RVT opB_reg_23_ ( .D(N92), .CLK(clk), .Q(opB[23]) );
  DFFX1_RVT opB_reg_22_ ( .D(N91), .CLK(clk), .Q(opB[22]) );
  DFFX1_RVT opB_reg_21_ ( .D(N90), .CLK(clk), .Q(opB[21]) );
  DFFX1_RVT opB_reg_20_ ( .D(N89), .CLK(clk), .Q(opB[20]) );
  DFFX1_RVT opB_reg_19_ ( .D(N88), .CLK(clk), .Q(opB[19]) );
  DFFX1_RVT opB_reg_18_ ( .D(N87), .CLK(clk), .Q(opB[18]) );
  DFFX1_RVT opB_reg_17_ ( .D(N86), .CLK(clk), .Q(opB[17]) );
  DFFX1_RVT opB_reg_16_ ( .D(N85), .CLK(clk), .Q(opB[16]) );
  DFFX1_RVT opB_reg_15_ ( .D(N84), .CLK(clk), .Q(opB[15]) );
  DFFX1_RVT opB_reg_14_ ( .D(N83), .CLK(clk), .Q(opB[14]) );
  DFFX1_RVT opB_reg_13_ ( .D(N82), .CLK(clk), .Q(opB[13]) );
  DFFX1_RVT opB_reg_12_ ( .D(N81), .CLK(clk), .Q(opB[12]) );
  DFFX1_RVT opB_reg_11_ ( .D(N80), .CLK(clk), .Q(opB[11]) );
  DFFX1_RVT opB_reg_10_ ( .D(N79), .CLK(clk), .Q(opB[10]) );
  DFFX1_RVT opB_reg_9_ ( .D(N78), .CLK(clk), .Q(opB[9]) );
  DFFX1_RVT opB_reg_8_ ( .D(N77), .CLK(clk), .Q(opB[8]) );
  DFFX1_RVT opB_reg_7_ ( .D(N76), .CLK(clk), .Q(opB[7]) );
  DFFX1_RVT opB_reg_6_ ( .D(N75), .CLK(clk), .Q(opB[6]) );
  DFFX1_RVT opB_reg_5_ ( .D(N74), .CLK(clk), .Q(opB[5]) );
  DFFX1_RVT opB_reg_4_ ( .D(N73), .CLK(clk), .Q(opB[4]) );
  DFFX1_RVT opB_reg_3_ ( .D(N72), .CLK(clk), .Q(opB[3]) );
  DFFX1_RVT opB_reg_2_ ( .D(N71), .CLK(clk), .Q(opB[2]) );
  DFFX1_RVT opB_reg_1_ ( .D(N70), .CLK(clk), .Q(opB[1]) );
  DFFX1_RVT opB_reg_0_ ( .D(N69), .CLK(clk), .Q(opB[0]) );
  NBUFFX2_RVT U99 ( .A(rstnPipe), .Y(n2) );
  NBUFFX2_RVT U100 ( .A(rstnPipe), .Y(n4) );
  NBUFFX2_RVT U101 ( .A(rstnPipe), .Y(n3) );
  NBUFFX2_RVT U102 ( .A(rstnPipe), .Y(n1) );
  NBUFFX2_RVT U103 ( .A(rstnPipe), .Y(n5) );
  NBUFFX2_RVT U104 ( .A(rstnPsum), .Y(n6) );
  NBUFFX2_RVT U105 ( .A(rstnPsum), .Y(n7) );
endmodule


module OSPEArray ( clk, rstnPipe, rstnPsum, ipA0, ipA1, ipA2, ipA3, ipB0, ipB1, 
        ipB2, ipB3, opC00, opC01, opC02, opC03, opC10, opC11, opC12, opC13, 
        opC20, opC21, opC22, opC23, opC30, opC31, opC32, opC33 );
  input [15:0] rstnPsum;
  input [31:0] ipA0;
  input [31:0] ipA1;
  input [31:0] ipA2;
  input [31:0] ipA3;
  input [31:0] ipB0;
  input [31:0] ipB1;
  input [31:0] ipB2;
  input [31:0] ipB3;
  output [31:0] opC00;
  output [31:0] opC01;
  output [31:0] opC02;
  output [31:0] opC03;
  output [31:0] opC10;
  output [31:0] opC11;
  output [31:0] opC12;
  output [31:0] opC13;
  output [31:0] opC20;
  output [31:0] opC21;
  output [31:0] opC22;
  output [31:0] opC23;
  output [31:0] opC30;
  output [31:0] opC31;
  output [31:0] opC32;
  output [31:0] opC33;
  input clk, rstnPipe;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317,
         N318, N319, N320, N321, N322, N323, n3, n4, n7, n8, n11, n12, n15,
         n16, n19, n20, n23, n24, n27, n28, n31, n32, n35, n36, n39, n40, n43,
         n44, n47, n48, n51, n52, n55, n56, n59, n60, n63, n64, n67, n68, n71,
         n72, n75, n76, n79, n80, n83, n84, n87, n88, n91, n92, n95, n96, n99,
         n100, n103, n104, n107, n108, n111, n112, n115, n116, n119, n120,
         n123, n124, n127, n128, n162, n164, n166, n168, n170, n172, n174,
         n176, n178, n180, n182, n184, n186, n188, n190, n192, n194, n196,
         n198, n200, n202, n204, n206, n208, n210, n212, n214, n216, n218,
         n220, n222, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256;
  wire   [31:0] ipA1_d1;
  wire   [31:0] ipB1_d1;
  wire   [31:0] ipA2_d2;
  wire   [31:0] ipB2_d2;
  wire   [31:0] ipA3_d3;
  wire   [31:0] ipB3_d3;
  wire   [31:0] opA00;
  wire   [31:0] opB00;
  wire   [31:0] opA01;
  wire   [31:0] opB01;
  wire   [31:0] opA02;
  wire   [31:0] opB02;
  wire   [31:0] opB03;
  wire   [31:0] opA10;
  wire   [31:0] opB10;
  wire   [31:0] opA11;
  wire   [31:0] opB11;
  wire   [31:0] opA12;
  wire   [31:0] opB12;
  wire   [31:0] opB13;
  wire   [31:0] opA20;
  wire   [31:0] opB20;
  wire   [31:0] opA21;
  wire   [31:0] opB21;
  wire   [31:0] opA22;
  wire   [31:0] opB22;
  wire   [31:0] opB23;
  wire   [31:0] opA30;
  wire   [31:0] opA31;
  wire   [31:0] opA32;

  SDFFX1_RVT ipA2_d2_reg_31_ ( .D(n397), .SI(1'b0), .SE(n384), .CLK(clk), .Q(
        ipA2_d2[31]) );
  SDFFX1_RVT ipA2_d2_reg_30_ ( .D(n407), .SI(1'b0), .SE(n383), .CLK(clk), .Q(
        ipA2_d2[30]) );
  SDFFX1_RVT ipA2_d2_reg_29_ ( .D(n402), .SI(1'b0), .SE(n382), .CLK(clk), .Q(
        ipA2_d2[29]) );
  SDFFX1_RVT ipA2_d2_reg_28_ ( .D(n404), .SI(1'b0), .SE(n381), .CLK(clk), .Q(
        ipA2_d2[28]) );
  SDFFX1_RVT ipA2_d2_reg_27_ ( .D(n403), .SI(1'b0), .SE(n380), .CLK(clk), .Q(
        ipA2_d2[27]) );
  SDFFX1_RVT ipA2_d2_reg_26_ ( .D(n402), .SI(1'b0), .SE(n379), .CLK(clk), .Q(
        ipA2_d2[26]) );
  SDFFX1_RVT ipA2_d2_reg_25_ ( .D(n404), .SI(1'b0), .SE(n378), .CLK(clk), .Q(
        ipA2_d2[25]) );
  SDFFX1_RVT ipA2_d2_reg_24_ ( .D(n403), .SI(1'b0), .SE(n377), .CLK(clk), .Q(
        ipA2_d2[24]) );
  SDFFX1_RVT ipA2_d2_reg_23_ ( .D(n402), .SI(1'b0), .SE(n376), .CLK(clk), .Q(
        ipA2_d2[23]) );
  SDFFX1_RVT ipA2_d2_reg_22_ ( .D(n404), .SI(1'b0), .SE(n375), .CLK(clk), .Q(
        ipA2_d2[22]) );
  SDFFX1_RVT ipA2_d2_reg_21_ ( .D(n403), .SI(1'b0), .SE(n374), .CLK(clk), .Q(
        ipA2_d2[21]) );
  SDFFX1_RVT ipA2_d2_reg_20_ ( .D(n402), .SI(1'b0), .SE(n373), .CLK(clk), .Q(
        ipA2_d2[20]) );
  SDFFX1_RVT ipA2_d2_reg_19_ ( .D(n404), .SI(1'b0), .SE(n372), .CLK(clk), .Q(
        ipA2_d2[19]) );
  SDFFX1_RVT ipA2_d2_reg_18_ ( .D(n403), .SI(1'b0), .SE(n371), .CLK(clk), .Q(
        ipA2_d2[18]) );
  SDFFX1_RVT ipA2_d2_reg_17_ ( .D(n402), .SI(1'b0), .SE(n370), .CLK(clk), .Q(
        ipA2_d2[17]) );
  SDFFX1_RVT ipA2_d2_reg_16_ ( .D(n404), .SI(1'b0), .SE(n369), .CLK(clk), .Q(
        ipA2_d2[16]) );
  SDFFX1_RVT ipA2_d2_reg_15_ ( .D(n403), .SI(1'b0), .SE(n368), .CLK(clk), .Q(
        ipA2_d2[15]) );
  SDFFX1_RVT ipA2_d2_reg_14_ ( .D(n402), .SI(1'b0), .SE(n367), .CLK(clk), .Q(
        ipA2_d2[14]) );
  SDFFX1_RVT ipA2_d2_reg_13_ ( .D(n404), .SI(1'b0), .SE(n366), .CLK(clk), .Q(
        ipA2_d2[13]) );
  SDFFX1_RVT ipA2_d2_reg_12_ ( .D(n403), .SI(1'b0), .SE(n365), .CLK(clk), .Q(
        ipA2_d2[12]) );
  SDFFX1_RVT ipA2_d2_reg_11_ ( .D(n402), .SI(1'b0), .SE(n364), .CLK(clk), .Q(
        ipA2_d2[11]) );
  SDFFX1_RVT ipA2_d2_reg_10_ ( .D(n404), .SI(1'b0), .SE(n363), .CLK(clk), .Q(
        ipA2_d2[10]) );
  SDFFX1_RVT ipA2_d2_reg_9_ ( .D(n403), .SI(1'b0), .SE(n362), .CLK(clk), .Q(
        ipA2_d2[9]) );
  SDFFX1_RVT ipA2_d2_reg_8_ ( .D(n402), .SI(1'b0), .SE(n361), .CLK(clk), .Q(
        ipA2_d2[8]) );
  SDFFX1_RVT ipA2_d2_reg_7_ ( .D(n404), .SI(1'b0), .SE(n360), .CLK(clk), .Q(
        ipA2_d2[7]) );
  SDFFX1_RVT ipA2_d2_reg_6_ ( .D(n403), .SI(1'b0), .SE(n359), .CLK(clk), .Q(
        ipA2_d2[6]) );
  SDFFX1_RVT ipA2_d2_reg_5_ ( .D(n402), .SI(1'b0), .SE(n358), .CLK(clk), .Q(
        ipA2_d2[5]) );
  SDFFX1_RVT ipA2_d2_reg_4_ ( .D(n404), .SI(1'b0), .SE(n357), .CLK(clk), .Q(
        ipA2_d2[4]) );
  SDFFX1_RVT ipA2_d2_reg_3_ ( .D(n403), .SI(1'b0), .SE(n356), .CLK(clk), .Q(
        ipA2_d2[3]) );
  SDFFX1_RVT ipA2_d2_reg_2_ ( .D(n402), .SI(1'b0), .SE(n355), .CLK(clk), .Q(
        ipA2_d2[2]) );
  SDFFX1_RVT ipA2_d2_reg_1_ ( .D(n404), .SI(1'b0), .SE(n354), .CLK(clk), .Q(
        ipA2_d2[1]) );
  SDFFX1_RVT ipA2_d2_reg_0_ ( .D(n403), .SI(1'b0), .SE(n353), .CLK(clk), .Q(
        ipA2_d2[0]) );
  SDFFX1_RVT ipB2_d2_reg_31_ ( .D(n402), .SI(1'b0), .SE(n320), .CLK(clk), .Q(
        ipB2_d2[31]) );
  SDFFX1_RVT ipB2_d2_reg_30_ ( .D(n406), .SI(1'b0), .SE(n319), .CLK(clk), .Q(
        ipB2_d2[30]) );
  SDFFX1_RVT ipB2_d2_reg_29_ ( .D(n405), .SI(1'b0), .SE(n318), .CLK(clk), .Q(
        ipB2_d2[29]) );
  SDFFX1_RVT ipB2_d2_reg_28_ ( .D(n407), .SI(1'b0), .SE(n317), .CLK(clk), .Q(
        ipB2_d2[28]) );
  SDFFX1_RVT ipB2_d2_reg_27_ ( .D(n406), .SI(1'b0), .SE(n316), .CLK(clk), .Q(
        ipB2_d2[27]) );
  SDFFX1_RVT ipB2_d2_reg_26_ ( .D(n405), .SI(1'b0), .SE(n315), .CLK(clk), .Q(
        ipB2_d2[26]) );
  SDFFX1_RVT ipB2_d2_reg_25_ ( .D(n407), .SI(1'b0), .SE(n314), .CLK(clk), .Q(
        ipB2_d2[25]) );
  SDFFX1_RVT ipB2_d2_reg_24_ ( .D(n406), .SI(1'b0), .SE(n313), .CLK(clk), .Q(
        ipB2_d2[24]) );
  SDFFX1_RVT ipB2_d2_reg_23_ ( .D(n405), .SI(1'b0), .SE(n312), .CLK(clk), .Q(
        ipB2_d2[23]) );
  SDFFX1_RVT ipB2_d2_reg_22_ ( .D(n407), .SI(1'b0), .SE(n311), .CLK(clk), .Q(
        ipB2_d2[22]) );
  SDFFX1_RVT ipB2_d2_reg_21_ ( .D(n406), .SI(1'b0), .SE(n310), .CLK(clk), .Q(
        ipB2_d2[21]) );
  SDFFX1_RVT ipB2_d2_reg_20_ ( .D(n405), .SI(1'b0), .SE(n309), .CLK(clk), .Q(
        ipB2_d2[20]) );
  SDFFX1_RVT ipB2_d2_reg_19_ ( .D(n407), .SI(1'b0), .SE(n308), .CLK(clk), .Q(
        ipB2_d2[19]) );
  SDFFX1_RVT ipB2_d2_reg_18_ ( .D(n406), .SI(1'b0), .SE(n307), .CLK(clk), .Q(
        ipB2_d2[18]) );
  SDFFX1_RVT ipB2_d2_reg_17_ ( .D(n405), .SI(1'b0), .SE(n306), .CLK(clk), .Q(
        ipB2_d2[17]) );
  SDFFX1_RVT ipB2_d2_reg_16_ ( .D(n407), .SI(1'b0), .SE(n305), .CLK(clk), .Q(
        ipB2_d2[16]) );
  SDFFX1_RVT ipB2_d2_reg_15_ ( .D(n406), .SI(1'b0), .SE(n304), .CLK(clk), .Q(
        ipB2_d2[15]) );
  SDFFX1_RVT ipB2_d2_reg_14_ ( .D(n405), .SI(1'b0), .SE(n303), .CLK(clk), .Q(
        ipB2_d2[14]) );
  SDFFX1_RVT ipB2_d2_reg_13_ ( .D(n407), .SI(1'b0), .SE(n302), .CLK(clk), .Q(
        ipB2_d2[13]) );
  SDFFX1_RVT ipB2_d2_reg_12_ ( .D(n406), .SI(1'b0), .SE(n301), .CLK(clk), .Q(
        ipB2_d2[12]) );
  SDFFX1_RVT ipB2_d2_reg_11_ ( .D(n405), .SI(1'b0), .SE(n300), .CLK(clk), .Q(
        ipB2_d2[11]) );
  SDFFX1_RVT ipB2_d2_reg_10_ ( .D(n406), .SI(1'b0), .SE(n299), .CLK(clk), .Q(
        ipB2_d2[10]) );
  SDFFX1_RVT ipB2_d2_reg_9_ ( .D(n405), .SI(1'b0), .SE(n298), .CLK(clk), .Q(
        ipB2_d2[9]) );
  SDFFX1_RVT ipB2_d2_reg_8_ ( .D(n407), .SI(1'b0), .SE(n297), .CLK(clk), .Q(
        ipB2_d2[8]) );
  SDFFX1_RVT ipB2_d2_reg_7_ ( .D(n406), .SI(1'b0), .SE(n296), .CLK(clk), .Q(
        ipB2_d2[7]) );
  SDFFX1_RVT ipB2_d2_reg_6_ ( .D(n405), .SI(1'b0), .SE(n295), .CLK(clk), .Q(
        ipB2_d2[6]) );
  SDFFX1_RVT ipB2_d2_reg_5_ ( .D(n407), .SI(1'b0), .SE(n294), .CLK(clk), .Q(
        ipB2_d2[5]) );
  SDFFX1_RVT ipB2_d2_reg_4_ ( .D(n406), .SI(1'b0), .SE(n293), .CLK(clk), .Q(
        ipB2_d2[4]) );
  SDFFX1_RVT ipB2_d2_reg_3_ ( .D(n405), .SI(1'b0), .SE(n292), .CLK(clk), .Q(
        ipB2_d2[3]) );
  SDFFX1_RVT ipB2_d2_reg_2_ ( .D(n407), .SI(1'b0), .SE(n291), .CLK(clk), .Q(
        ipB2_d2[2]) );
  SDFFX1_RVT ipB2_d2_reg_1_ ( .D(n406), .SI(1'b0), .SE(n290), .CLK(clk), .Q(
        ipB2_d2[1]) );
  SDFFX1_RVT ipB2_d2_reg_0_ ( .D(n405), .SI(1'b0), .SE(n289), .CLK(clk), .Q(
        ipB2_d2[0]) );
  SDFFX1_RVT ipA3_d2_reg_31_ ( .D(n407), .SI(1'b0), .SE(n256), .CLK(clk), .QN(
        n224) );
  SDFFX1_RVT ipA3_d2_reg_30_ ( .D(n406), .SI(1'b0), .SE(n255), .CLK(clk), .QN(
        n222) );
  SDFFX1_RVT ipA3_d2_reg_29_ ( .D(n405), .SI(1'b0), .SE(n254), .CLK(clk), .QN(
        n220) );
  SDFFX1_RVT ipA3_d2_reg_28_ ( .D(n407), .SI(1'b0), .SE(n253), .CLK(clk), .QN(
        n218) );
  SDFFX1_RVT ipA3_d2_reg_27_ ( .D(n406), .SI(1'b0), .SE(n252), .CLK(clk), .QN(
        n216) );
  SDFFX1_RVT ipA3_d2_reg_26_ ( .D(n405), .SI(1'b0), .SE(n251), .CLK(clk), .QN(
        n214) );
  SDFFX1_RVT ipA3_d2_reg_25_ ( .D(n407), .SI(1'b0), .SE(n250), .CLK(clk), .QN(
        n212) );
  SDFFX1_RVT ipA3_d2_reg_24_ ( .D(n406), .SI(1'b0), .SE(n249), .CLK(clk), .QN(
        n210) );
  SDFFX1_RVT ipA3_d2_reg_23_ ( .D(n405), .SI(1'b0), .SE(n248), .CLK(clk), .QN(
        n208) );
  SDFFX1_RVT ipA3_d2_reg_22_ ( .D(n407), .SI(1'b0), .SE(n247), .CLK(clk), .QN(
        n206) );
  SDFFX1_RVT ipA3_d2_reg_21_ ( .D(n406), .SI(1'b0), .SE(n246), .CLK(clk), .QN(
        n204) );
  SDFFX1_RVT ipA3_d2_reg_20_ ( .D(n405), .SI(1'b0), .SE(n245), .CLK(clk), .QN(
        n202) );
  SDFFX1_RVT ipA3_d2_reg_19_ ( .D(n407), .SI(1'b0), .SE(n244), .CLK(clk), .QN(
        n200) );
  SDFFX1_RVT ipA3_d2_reg_18_ ( .D(n406), .SI(1'b0), .SE(n243), .CLK(clk), .QN(
        n198) );
  SDFFX1_RVT ipA3_d2_reg_17_ ( .D(n405), .SI(1'b0), .SE(n242), .CLK(clk), .QN(
        n196) );
  SDFFX1_RVT ipA3_d2_reg_16_ ( .D(n407), .SI(1'b0), .SE(n241), .CLK(clk), .QN(
        n194) );
  SDFFX1_RVT ipA3_d2_reg_15_ ( .D(n406), .SI(1'b0), .SE(n240), .CLK(clk), .QN(
        n192) );
  SDFFX1_RVT ipA3_d2_reg_14_ ( .D(n405), .SI(1'b0), .SE(n239), .CLK(clk), .QN(
        n190) );
  SDFFX1_RVT ipA3_d2_reg_13_ ( .D(n409), .SI(1'b0), .SE(n238), .CLK(clk), .QN(
        n188) );
  SDFFX1_RVT ipA3_d2_reg_12_ ( .D(n410), .SI(1'b0), .SE(n237), .CLK(clk), .QN(
        n186) );
  SDFFX1_RVT ipA3_d2_reg_11_ ( .D(n409), .SI(1'b0), .SE(n236), .CLK(clk), .QN(
        n184) );
  SDFFX1_RVT ipA3_d2_reg_10_ ( .D(n410), .SI(1'b0), .SE(n235), .CLK(clk), .QN(
        n182) );
  SDFFX1_RVT ipA3_d2_reg_9_ ( .D(n409), .SI(1'b0), .SE(n234), .CLK(clk), .QN(
        n180) );
  SDFFX1_RVT ipA3_d2_reg_8_ ( .D(n410), .SI(1'b0), .SE(n233), .CLK(clk), .QN(
        n178) );
  SDFFX1_RVT ipA3_d2_reg_7_ ( .D(n409), .SI(1'b0), .SE(n232), .CLK(clk), .QN(
        n176) );
  SDFFX1_RVT ipA3_d2_reg_6_ ( .D(n410), .SI(1'b0), .SE(n231), .CLK(clk), .QN(
        n174) );
  SDFFX1_RVT ipA3_d2_reg_5_ ( .D(n409), .SI(1'b0), .SE(n230), .CLK(clk), .QN(
        n172) );
  SDFFX1_RVT ipA3_d2_reg_4_ ( .D(n410), .SI(1'b0), .SE(n229), .CLK(clk), .QN(
        n170) );
  SDFFX1_RVT ipA3_d2_reg_3_ ( .D(n409), .SI(1'b0), .SE(n228), .CLK(clk), .QN(
        n168) );
  SDFFX1_RVT ipA3_d2_reg_2_ ( .D(n410), .SI(1'b0), .SE(n227), .CLK(clk), .QN(
        n166) );
  SDFFX1_RVT ipA3_d2_reg_1_ ( .D(n409), .SI(1'b0), .SE(n226), .CLK(clk), .QN(
        n164) );
  SDFFX1_RVT ipA3_d2_reg_0_ ( .D(n410), .SI(1'b0), .SE(n225), .CLK(clk), .QN(
        n162) );
  SDFFX1_RVT ipA3_d3_reg_31_ ( .D(n408), .SI(1'b0), .SE(n224), .CLK(clk), .Q(
        ipA3_d3[31]) );
  SDFFX1_RVT ipA3_d3_reg_30_ ( .D(n408), .SI(1'b0), .SE(n222), .CLK(clk), .Q(
        ipA3_d3[30]) );
  SDFFX1_RVT ipA3_d3_reg_29_ ( .D(n408), .SI(1'b0), .SE(n220), .CLK(clk), .Q(
        ipA3_d3[29]) );
  SDFFX1_RVT ipA3_d3_reg_28_ ( .D(n408), .SI(1'b0), .SE(n218), .CLK(clk), .Q(
        ipA3_d3[28]) );
  SDFFX1_RVT ipA3_d3_reg_27_ ( .D(n408), .SI(1'b0), .SE(n216), .CLK(clk), .Q(
        ipA3_d3[27]) );
  SDFFX1_RVT ipA3_d3_reg_26_ ( .D(n408), .SI(1'b0), .SE(n214), .CLK(clk), .Q(
        ipA3_d3[26]) );
  SDFFX1_RVT ipA3_d3_reg_25_ ( .D(n408), .SI(1'b0), .SE(n212), .CLK(clk), .Q(
        ipA3_d3[25]) );
  SDFFX1_RVT ipA3_d3_reg_24_ ( .D(n408), .SI(1'b0), .SE(n210), .CLK(clk), .Q(
        ipA3_d3[24]) );
  SDFFX1_RVT ipA3_d3_reg_23_ ( .D(n401), .SI(1'b0), .SE(n208), .CLK(clk), .Q(
        ipA3_d3[23]) );
  SDFFX1_RVT ipA3_d3_reg_22_ ( .D(n398), .SI(1'b0), .SE(n206), .CLK(clk), .Q(
        ipA3_d3[22]) );
  SDFFX1_RVT ipA3_d3_reg_21_ ( .D(n397), .SI(1'b0), .SE(n204), .CLK(clk), .Q(
        ipA3_d3[21]) );
  SDFFX1_RVT ipA3_d3_reg_20_ ( .D(n403), .SI(1'b0), .SE(n202), .CLK(clk), .Q(
        ipA3_d3[20]) );
  SDFFX1_RVT ipA3_d3_reg_19_ ( .D(n398), .SI(1'b0), .SE(n200), .CLK(clk), .Q(
        ipA3_d3[19]) );
  SDFFX1_RVT ipA3_d3_reg_18_ ( .D(n397), .SI(1'b0), .SE(n198), .CLK(clk), .Q(
        ipA3_d3[18]) );
  SDFFX1_RVT ipA3_d3_reg_17_ ( .D(n398), .SI(1'b0), .SE(n196), .CLK(clk), .Q(
        ipA3_d3[17]) );
  SDFFX1_RVT ipA3_d3_reg_16_ ( .D(n397), .SI(1'b0), .SE(n194), .CLK(clk), .Q(
        ipA3_d3[16]) );
  SDFFX1_RVT ipA3_d3_reg_15_ ( .D(n398), .SI(1'b0), .SE(n192), .CLK(clk), .Q(
        ipA3_d3[15]) );
  SDFFX1_RVT ipA3_d3_reg_14_ ( .D(n397), .SI(1'b0), .SE(n190), .CLK(clk), .Q(
        ipA3_d3[14]) );
  SDFFX1_RVT ipA3_d3_reg_13_ ( .D(n398), .SI(1'b0), .SE(n188), .CLK(clk), .Q(
        ipA3_d3[13]) );
  SDFFX1_RVT ipA3_d3_reg_12_ ( .D(n397), .SI(1'b0), .SE(n186), .CLK(clk), .Q(
        ipA3_d3[12]) );
  SDFFX1_RVT ipA3_d3_reg_11_ ( .D(n398), .SI(1'b0), .SE(n184), .CLK(clk), .Q(
        ipA3_d3[11]) );
  SDFFX1_RVT ipA3_d3_reg_10_ ( .D(n397), .SI(1'b0), .SE(n182), .CLK(clk), .Q(
        ipA3_d3[10]) );
  SDFFX1_RVT ipA3_d3_reg_9_ ( .D(n398), .SI(1'b0), .SE(n180), .CLK(clk), .Q(
        ipA3_d3[9]) );
  SDFFX1_RVT ipA3_d3_reg_8_ ( .D(n397), .SI(1'b0), .SE(n178), .CLK(clk), .Q(
        ipA3_d3[8]) );
  SDFFX1_RVT ipA3_d3_reg_7_ ( .D(n398), .SI(1'b0), .SE(n176), .CLK(clk), .Q(
        ipA3_d3[7]) );
  SDFFX1_RVT ipA3_d3_reg_6_ ( .D(n397), .SI(1'b0), .SE(n174), .CLK(clk), .Q(
        ipA3_d3[6]) );
  SDFFX1_RVT ipA3_d3_reg_5_ ( .D(n398), .SI(1'b0), .SE(n172), .CLK(clk), .Q(
        ipA3_d3[5]) );
  SDFFX1_RVT ipA3_d3_reg_4_ ( .D(n397), .SI(1'b0), .SE(n170), .CLK(clk), .Q(
        ipA3_d3[4]) );
  SDFFX1_RVT ipA3_d3_reg_3_ ( .D(n398), .SI(1'b0), .SE(n168), .CLK(clk), .Q(
        ipA3_d3[3]) );
  SDFFX1_RVT ipA3_d3_reg_2_ ( .D(n400), .SI(1'b0), .SE(n166), .CLK(clk), .Q(
        ipA3_d3[2]) );
  SDFFX1_RVT ipA3_d3_reg_1_ ( .D(n399), .SI(1'b0), .SE(n164), .CLK(clk), .Q(
        ipA3_d3[1]) );
  SDFFX1_RVT ipA3_d3_reg_0_ ( .D(n401), .SI(1'b0), .SE(n162), .CLK(clk), .Q(
        ipA3_d3[0]) );
  SDFFX1_RVT ipB3_d2_reg_31_ ( .D(n400), .SI(1'b0), .SE(n128), .CLK(clk), .QN(
        n127) );
  SDFFX1_RVT ipB3_d3_reg_31_ ( .D(n399), .SI(1'b0), .SE(n127), .CLK(clk), .Q(
        ipB3_d3[31]) );
  SDFFX1_RVT ipB3_d2_reg_30_ ( .D(n401), .SI(1'b0), .SE(n124), .CLK(clk), .QN(
        n123) );
  SDFFX1_RVT ipB3_d3_reg_30_ ( .D(n400), .SI(1'b0), .SE(n123), .CLK(clk), .Q(
        ipB3_d3[30]) );
  SDFFX1_RVT ipB3_d2_reg_29_ ( .D(n399), .SI(1'b0), .SE(n120), .CLK(clk), .QN(
        n119) );
  SDFFX1_RVT ipB3_d3_reg_29_ ( .D(n401), .SI(1'b0), .SE(n119), .CLK(clk), .Q(
        ipB3_d3[29]) );
  SDFFX1_RVT ipB3_d2_reg_28_ ( .D(n400), .SI(1'b0), .SE(n116), .CLK(clk), .QN(
        n115) );
  SDFFX1_RVT ipB3_d3_reg_28_ ( .D(n399), .SI(1'b0), .SE(n115), .CLK(clk), .Q(
        ipB3_d3[28]) );
  SDFFX1_RVT ipB3_d2_reg_27_ ( .D(n401), .SI(1'b0), .SE(n112), .CLK(clk), .QN(
        n111) );
  SDFFX1_RVT ipB3_d3_reg_27_ ( .D(n400), .SI(1'b0), .SE(n111), .CLK(clk), .Q(
        ipB3_d3[27]) );
  SDFFX1_RVT ipB3_d2_reg_26_ ( .D(n399), .SI(1'b0), .SE(n108), .CLK(clk), .QN(
        n107) );
  SDFFX1_RVT ipB3_d3_reg_26_ ( .D(n401), .SI(1'b0), .SE(n107), .CLK(clk), .Q(
        ipB3_d3[26]) );
  SDFFX1_RVT ipB3_d2_reg_25_ ( .D(n400), .SI(1'b0), .SE(n104), .CLK(clk), .QN(
        n103) );
  SDFFX1_RVT ipB3_d3_reg_25_ ( .D(n399), .SI(1'b0), .SE(n103), .CLK(clk), .Q(
        ipB3_d3[25]) );
  SDFFX1_RVT ipB3_d2_reg_24_ ( .D(n401), .SI(1'b0), .SE(n100), .CLK(clk), .QN(
        n99) );
  SDFFX1_RVT ipB3_d3_reg_24_ ( .D(n400), .SI(1'b0), .SE(n99), .CLK(clk), .Q(
        ipB3_d3[24]) );
  SDFFX1_RVT ipB3_d2_reg_23_ ( .D(n399), .SI(1'b0), .SE(n96), .CLK(clk), .QN(
        n95) );
  SDFFX1_RVT ipB3_d3_reg_23_ ( .D(n401), .SI(1'b0), .SE(n95), .CLK(clk), .Q(
        ipB3_d3[23]) );
  SDFFX1_RVT ipB3_d2_reg_22_ ( .D(n400), .SI(1'b0), .SE(n92), .CLK(clk), .QN(
        n91) );
  SDFFX1_RVT ipB3_d3_reg_22_ ( .D(n399), .SI(1'b0), .SE(n91), .CLK(clk), .Q(
        ipB3_d3[22]) );
  SDFFX1_RVT ipB3_d2_reg_21_ ( .D(n400), .SI(1'b0), .SE(n88), .CLK(clk), .QN(
        n87) );
  SDFFX1_RVT ipB3_d3_reg_21_ ( .D(n399), .SI(1'b0), .SE(n87), .CLK(clk), .Q(
        ipB3_d3[21]) );
  SDFFX1_RVT ipB3_d2_reg_20_ ( .D(n401), .SI(1'b0), .SE(n84), .CLK(clk), .QN(
        n83) );
  SDFFX1_RVT ipB3_d3_reg_20_ ( .D(n400), .SI(1'b0), .SE(n83), .CLK(clk), .Q(
        ipB3_d3[20]) );
  SDFFX1_RVT ipB3_d2_reg_19_ ( .D(n399), .SI(1'b0), .SE(n80), .CLK(clk), .QN(
        n79) );
  SDFFX1_RVT ipB3_d3_reg_19_ ( .D(n401), .SI(1'b0), .SE(n79), .CLK(clk), .Q(
        ipB3_d3[19]) );
  SDFFX1_RVT ipB3_d2_reg_18_ ( .D(n400), .SI(1'b0), .SE(n76), .CLK(clk), .QN(
        n75) );
  SDFFX1_RVT ipB3_d3_reg_18_ ( .D(n399), .SI(1'b0), .SE(n75), .CLK(clk), .Q(
        ipB3_d3[18]) );
  SDFFX1_RVT ipB3_d2_reg_17_ ( .D(n401), .SI(1'b0), .SE(n72), .CLK(clk), .QN(
        n71) );
  SDFFX1_RVT ipB3_d3_reg_17_ ( .D(n400), .SI(1'b0), .SE(n71), .CLK(clk), .Q(
        ipB3_d3[17]) );
  SDFFX1_RVT ipB3_d2_reg_16_ ( .D(n399), .SI(1'b0), .SE(n68), .CLK(clk), .QN(
        n67) );
  SDFFX1_RVT ipB3_d3_reg_16_ ( .D(n401), .SI(1'b0), .SE(n67), .CLK(clk), .Q(
        ipB3_d3[16]) );
  SDFFX1_RVT ipB3_d2_reg_15_ ( .D(n400), .SI(1'b0), .SE(n64), .CLK(clk), .QN(
        n63) );
  SDFFX1_RVT ipB3_d3_reg_15_ ( .D(n399), .SI(1'b0), .SE(n63), .CLK(clk), .Q(
        ipB3_d3[15]) );
  SDFFX1_RVT ipB3_d2_reg_14_ ( .D(n401), .SI(1'b0), .SE(n60), .CLK(clk), .QN(
        n59) );
  SDFFX1_RVT ipB3_d3_reg_14_ ( .D(n400), .SI(1'b0), .SE(n59), .CLK(clk), .Q(
        ipB3_d3[14]) );
  SDFFX1_RVT ipB3_d2_reg_13_ ( .D(n399), .SI(1'b0), .SE(n56), .CLK(clk), .QN(
        n55) );
  SDFFX1_RVT ipB3_d3_reg_13_ ( .D(n401), .SI(1'b0), .SE(n55), .CLK(clk), .Q(
        ipB3_d3[13]) );
  SDFFX1_RVT ipB3_d2_reg_12_ ( .D(n400), .SI(1'b0), .SE(n52), .CLK(clk), .QN(
        n51) );
  SDFFX1_RVT ipB3_d3_reg_12_ ( .D(n399), .SI(1'b0), .SE(n51), .CLK(clk), .Q(
        ipB3_d3[12]) );
  SDFFX1_RVT ipB3_d2_reg_11_ ( .D(n401), .SI(1'b0), .SE(n48), .CLK(clk), .QN(
        n47) );
  SDFFX1_RVT ipB3_d3_reg_11_ ( .D(n400), .SI(1'b0), .SE(n47), .CLK(clk), .Q(
        ipB3_d3[11]) );
  SDFFX1_RVT ipB3_d2_reg_10_ ( .D(n399), .SI(1'b0), .SE(n44), .CLK(clk), .QN(
        n43) );
  SDFFX1_RVT ipB3_d3_reg_10_ ( .D(n401), .SI(1'b0), .SE(n43), .CLK(clk), .Q(
        ipB3_d3[10]) );
  SDFFX1_RVT ipB3_d2_reg_9_ ( .D(n400), .SI(1'b0), .SE(n40), .CLK(clk), .QN(
        n39) );
  SDFFX1_RVT ipB3_d3_reg_9_ ( .D(n399), .SI(1'b0), .SE(n39), .CLK(clk), .Q(
        ipB3_d3[9]) );
  SDFFX1_RVT ipB3_d2_reg_8_ ( .D(n403), .SI(1'b0), .SE(n36), .CLK(clk), .QN(
        n35) );
  SDFFX1_RVT ipB3_d3_reg_8_ ( .D(n402), .SI(1'b0), .SE(n35), .CLK(clk), .Q(
        ipB3_d3[8]) );
  SDFFX1_RVT ipB3_d2_reg_7_ ( .D(n404), .SI(1'b0), .SE(n32), .CLK(clk), .QN(
        n31) );
  SDFFX1_RVT ipB3_d3_reg_7_ ( .D(n403), .SI(1'b0), .SE(n31), .CLK(clk), .Q(
        ipB3_d3[7]) );
  SDFFX1_RVT ipB3_d2_reg_6_ ( .D(n402), .SI(1'b0), .SE(n28), .CLK(clk), .QN(
        n27) );
  SDFFX1_RVT ipB3_d3_reg_6_ ( .D(n404), .SI(1'b0), .SE(n27), .CLK(clk), .Q(
        ipB3_d3[6]) );
  SDFFX1_RVT ipB3_d2_reg_5_ ( .D(n403), .SI(1'b0), .SE(n24), .CLK(clk), .QN(
        n23) );
  SDFFX1_RVT ipB3_d3_reg_5_ ( .D(n402), .SI(1'b0), .SE(n23), .CLK(clk), .Q(
        ipB3_d3[5]) );
  SDFFX1_RVT ipB3_d2_reg_4_ ( .D(n404), .SI(1'b0), .SE(n20), .CLK(clk), .QN(
        n19) );
  SDFFX1_RVT ipB3_d3_reg_4_ ( .D(n403), .SI(1'b0), .SE(n19), .CLK(clk), .Q(
        ipB3_d3[4]) );
  SDFFX1_RVT ipB3_d2_reg_3_ ( .D(n402), .SI(1'b0), .SE(n16), .CLK(clk), .QN(
        n15) );
  SDFFX1_RVT ipB3_d3_reg_3_ ( .D(n404), .SI(1'b0), .SE(n15), .CLK(clk), .Q(
        ipB3_d3[3]) );
  SDFFX1_RVT ipB3_d2_reg_2_ ( .D(n403), .SI(1'b0), .SE(n12), .CLK(clk), .QN(
        n11) );
  SDFFX1_RVT ipB3_d3_reg_2_ ( .D(n402), .SI(1'b0), .SE(n11), .CLK(clk), .Q(
        ipB3_d3[2]) );
  SDFFX1_RVT ipB3_d2_reg_1_ ( .D(n404), .SI(1'b0), .SE(n8), .CLK(clk), .QN(n7)
         );
  SDFFX1_RVT ipB3_d3_reg_1_ ( .D(n403), .SI(1'b0), .SE(n7), .CLK(clk), .Q(
        ipB3_d3[1]) );
  SDFFX1_RVT ipB3_d2_reg_0_ ( .D(n402), .SI(1'b0), .SE(n4), .CLK(clk), .QN(n3)
         );
  SDFFX1_RVT ipB3_d3_reg_0_ ( .D(n404), .SI(1'b0), .SE(n3), .CLK(clk), .Q(
        ipB3_d3[0]) );
  AND2X1_RVT U195 ( .A1(n387), .A2(ipA2[31]), .Y(N99) );
  AND2X1_RVT U196 ( .A1(ipA2[30]), .A2(n386), .Y(N98) );
  AND2X1_RVT U197 ( .A1(ipA2[29]), .A2(n413), .Y(N97) );
  AND2X1_RVT U198 ( .A1(ipA2[28]), .A2(n391), .Y(N96) );
  AND2X1_RVT U199 ( .A1(ipA2[27]), .A2(n392), .Y(N95) );
  AND2X1_RVT U200 ( .A1(ipA2[26]), .A2(n414), .Y(N94) );
  AND2X1_RVT U201 ( .A1(ipA2[25]), .A2(n391), .Y(N93) );
  AND2X1_RVT U202 ( .A1(ipA2[24]), .A2(n392), .Y(N92) );
  AND2X1_RVT U203 ( .A1(ipA2[23]), .A2(n410), .Y(N91) );
  AND2X1_RVT U204 ( .A1(ipA2[22]), .A2(n391), .Y(N90) );
  AND2X1_RVT U205 ( .A1(ipA1[5]), .A2(n392), .Y(N9) );
  AND2X1_RVT U206 ( .A1(ipA2[21]), .A2(n413), .Y(N89) );
  AND2X1_RVT U207 ( .A1(ipA2[20]), .A2(n391), .Y(N88) );
  AND2X1_RVT U208 ( .A1(ipA2[19]), .A2(n392), .Y(N87) );
  AND2X1_RVT U209 ( .A1(ipA2[18]), .A2(n414), .Y(N86) );
  AND2X1_RVT U210 ( .A1(ipA2[17]), .A2(n388), .Y(N85) );
  AND2X1_RVT U211 ( .A1(ipA2[16]), .A2(n389), .Y(N84) );
  AND2X1_RVT U212 ( .A1(ipA2[15]), .A2(n390), .Y(N83) );
  AND2X1_RVT U213 ( .A1(ipA2[14]), .A2(n388), .Y(N82) );
  AND2X1_RVT U214 ( .A1(ipA2[13]), .A2(n389), .Y(N81) );
  AND2X1_RVT U215 ( .A1(ipA2[12]), .A2(n390), .Y(N80) );
  AND2X1_RVT U216 ( .A1(ipA1[4]), .A2(n388), .Y(N8) );
  AND2X1_RVT U217 ( .A1(ipA2[11]), .A2(n389), .Y(N79) );
  AND2X1_RVT U218 ( .A1(ipA2[10]), .A2(n390), .Y(N78) );
  AND2X1_RVT U219 ( .A1(ipA2[9]), .A2(n388), .Y(N77) );
  AND2X1_RVT U220 ( .A1(ipA2[8]), .A2(n389), .Y(N76) );
  AND2X1_RVT U221 ( .A1(ipA2[7]), .A2(n390), .Y(N75) );
  AND2X1_RVT U222 ( .A1(ipA2[6]), .A2(n388), .Y(N74) );
  AND2X1_RVT U223 ( .A1(ipA2[5]), .A2(n389), .Y(N73) );
  AND2X1_RVT U224 ( .A1(ipA2[4]), .A2(n390), .Y(N72) );
  AND2X1_RVT U225 ( .A1(ipA2[3]), .A2(n388), .Y(N71) );
  AND2X1_RVT U226 ( .A1(ipA2[2]), .A2(n389), .Y(N70) );
  AND2X1_RVT U227 ( .A1(ipA1[3]), .A2(n390), .Y(N7) );
  AND2X1_RVT U228 ( .A1(ipA2[1]), .A2(n388), .Y(N69) );
  AND2X1_RVT U229 ( .A1(ipA2[0]), .A2(n389), .Y(N68) );
  AND2X1_RVT U230 ( .A1(ipB1[31]), .A2(n390), .Y(N67) );
  AND2X1_RVT U231 ( .A1(ipB1[30]), .A2(n388), .Y(N66) );
  AND2X1_RVT U232 ( .A1(ipB1[29]), .A2(n389), .Y(N65) );
  AND2X1_RVT U233 ( .A1(ipB1[28]), .A2(n390), .Y(N64) );
  AND2X1_RVT U234 ( .A1(ipB1[27]), .A2(n388), .Y(N63) );
  AND2X1_RVT U235 ( .A1(ipB1[26]), .A2(n389), .Y(N62) );
  AND2X1_RVT U236 ( .A1(ipB1[25]), .A2(n390), .Y(N61) );
  AND2X1_RVT U237 ( .A1(ipB1[24]), .A2(n388), .Y(N60) );
  AND2X1_RVT U238 ( .A1(ipA1[2]), .A2(n389), .Y(N6) );
  AND2X1_RVT U239 ( .A1(ipB1[23]), .A2(n390), .Y(N59) );
  AND2X1_RVT U240 ( .A1(ipB1[22]), .A2(n389), .Y(N58) );
  AND2X1_RVT U241 ( .A1(ipB1[21]), .A2(n390), .Y(N57) );
  AND2X1_RVT U242 ( .A1(ipB1[20]), .A2(n388), .Y(N56) );
  AND2X1_RVT U243 ( .A1(ipB1[19]), .A2(n389), .Y(N55) );
  AND2X1_RVT U244 ( .A1(ipB1[18]), .A2(n390), .Y(N54) );
  AND2X1_RVT U245 ( .A1(ipB1[17]), .A2(n388), .Y(N53) );
  AND2X1_RVT U246 ( .A1(ipB1[16]), .A2(n389), .Y(N52) );
  AND2X1_RVT U247 ( .A1(ipB1[15]), .A2(n390), .Y(N51) );
  AND2X1_RVT U248 ( .A1(ipB1[14]), .A2(n388), .Y(N50) );
  AND2X1_RVT U249 ( .A1(ipA1[1]), .A2(n389), .Y(N5) );
  AND2X1_RVT U250 ( .A1(ipB1[13]), .A2(n390), .Y(N49) );
  AND2X1_RVT U251 ( .A1(ipB1[12]), .A2(n388), .Y(N48) );
  AND2X1_RVT U252 ( .A1(ipB1[11]), .A2(n389), .Y(N47) );
  AND2X1_RVT U253 ( .A1(ipB1[10]), .A2(n390), .Y(N46) );
  AND2X1_RVT U254 ( .A1(ipB1[9]), .A2(n386), .Y(N45) );
  AND2X1_RVT U255 ( .A1(ipB1[8]), .A2(n387), .Y(N44) );
  AND2X1_RVT U256 ( .A1(ipB1[7]), .A2(n386), .Y(N43) );
  AND2X1_RVT U257 ( .A1(ipB1[6]), .A2(n387), .Y(N42) );
  AND2X1_RVT U258 ( .A1(ipB1[5]), .A2(n386), .Y(N41) );
  AND2X1_RVT U259 ( .A1(ipB1[4]), .A2(n387), .Y(N40) );
  AND2X1_RVT U260 ( .A1(ipA1[0]), .A2(n386), .Y(N4) );
  AND2X1_RVT U261 ( .A1(ipB1[3]), .A2(n387), .Y(N39) );
  AND2X1_RVT U262 ( .A1(ipB1[2]), .A2(n386), .Y(N38) );
  AND2X1_RVT U263 ( .A1(ipB1[1]), .A2(n387), .Y(N37) );
  AND2X1_RVT U264 ( .A1(ipB1[0]), .A2(n386), .Y(N36) );
  AND2X1_RVT U265 ( .A1(ipA1[31]), .A2(n387), .Y(N35) );
  AND2X1_RVT U266 ( .A1(ipA1[30]), .A2(n386), .Y(N34) );
  AND2X1_RVT U267 ( .A1(ipA1[29]), .A2(n387), .Y(N33) );
  AND2X1_RVT U268 ( .A1(ipB3[31]), .A2(n386), .Y(N323) );
  AND2X1_RVT U269 ( .A1(ipB3[30]), .A2(n387), .Y(N322) );
  AND2X1_RVT U270 ( .A1(ipB3[29]), .A2(n386), .Y(N321) );
  AND2X1_RVT U271 ( .A1(ipB3[28]), .A2(n387), .Y(N320) );
  AND2X1_RVT U272 ( .A1(ipA1[28]), .A2(n386), .Y(N32) );
  AND2X1_RVT U273 ( .A1(ipB3[27]), .A2(n387), .Y(N319) );
  AND2X1_RVT U274 ( .A1(ipB3[26]), .A2(n386), .Y(N318) );
  AND2X1_RVT U275 ( .A1(ipB3[25]), .A2(n387), .Y(N317) );
  AND2X1_RVT U276 ( .A1(ipB3[24]), .A2(n386), .Y(N316) );
  AND2X1_RVT U277 ( .A1(ipB3[23]), .A2(n387), .Y(N315) );
  AND2X1_RVT U278 ( .A1(ipB3[22]), .A2(n386), .Y(N314) );
  AND2X1_RVT U279 ( .A1(ipB3[21]), .A2(n387), .Y(N313) );
  AND2X1_RVT U280 ( .A1(ipB3[20]), .A2(n386), .Y(N312) );
  AND2X1_RVT U281 ( .A1(ipB3[19]), .A2(n387), .Y(N311) );
  AND2X1_RVT U282 ( .A1(ipB3[18]), .A2(n388), .Y(N310) );
  AND2X1_RVT U283 ( .A1(ipA1[27]), .A2(n396), .Y(N31) );
  AND2X1_RVT U284 ( .A1(ipB3[17]), .A2(n396), .Y(N309) );
  AND2X1_RVT U285 ( .A1(ipB3[16]), .A2(n396), .Y(N308) );
  AND2X1_RVT U286 ( .A1(ipB3[15]), .A2(n396), .Y(N307) );
  AND2X1_RVT U287 ( .A1(ipB3[14]), .A2(n396), .Y(N306) );
  AND2X1_RVT U288 ( .A1(ipB3[13]), .A2(n396), .Y(N305) );
  AND2X1_RVT U289 ( .A1(ipB3[12]), .A2(n396), .Y(N304) );
  AND2X1_RVT U290 ( .A1(ipB3[11]), .A2(n396), .Y(N303) );
  AND2X1_RVT U291 ( .A1(ipB3[10]), .A2(n396), .Y(N302) );
  AND2X1_RVT U292 ( .A1(ipB3[9]), .A2(n396), .Y(N301) );
  AND2X1_RVT U293 ( .A1(ipB3[8]), .A2(n396), .Y(N300) );
  AND2X1_RVT U294 ( .A1(ipA1[26]), .A2(n396), .Y(N30) );
  AND2X1_RVT U295 ( .A1(ipB3[7]), .A2(n396), .Y(N299) );
  AND2X1_RVT U296 ( .A1(ipB3[6]), .A2(n396), .Y(N298) );
  AND2X1_RVT U297 ( .A1(ipB3[5]), .A2(n396), .Y(N297) );
  AND2X1_RVT U298 ( .A1(ipB3[4]), .A2(n398), .Y(N296) );
  AND2X1_RVT U299 ( .A1(ipB3[3]), .A2(n397), .Y(N295) );
  AND2X1_RVT U300 ( .A1(ipB3[2]), .A2(n398), .Y(N294) );
  AND2X1_RVT U301 ( .A1(ipB3[1]), .A2(n397), .Y(N293) );
  AND2X1_RVT U302 ( .A1(ipB3[0]), .A2(n398), .Y(N292) );
  AND2X1_RVT U303 ( .A1(ipA1[25]), .A2(n397), .Y(N29) );
  AND2X1_RVT U304 ( .A1(ipA1[24]), .A2(n398), .Y(N28) );
  AND2X1_RVT U305 ( .A1(ipA1[23]), .A2(n397), .Y(N27) );
  AND2X1_RVT U306 ( .A1(ipA1[22]), .A2(n398), .Y(N26) );
  AND2X1_RVT U307 ( .A1(ipA1[21]), .A2(n397), .Y(N25) );
  AND2X1_RVT U308 ( .A1(ipA1[20]), .A2(n398), .Y(N24) );
  AND2X1_RVT U309 ( .A1(ipA1[19]), .A2(n397), .Y(N23) );
  AND2X1_RVT U310 ( .A1(ipA3[31]), .A2(n393), .Y(N227) );
  AND2X1_RVT U311 ( .A1(ipA3[30]), .A2(n394), .Y(N226) );
  AND2X1_RVT U312 ( .A1(ipA3[29]), .A2(n395), .Y(N225) );
  AND2X1_RVT U313 ( .A1(ipA3[28]), .A2(n393), .Y(N224) );
  AND2X1_RVT U314 ( .A1(ipA3[27]), .A2(n394), .Y(N223) );
  AND2X1_RVT U315 ( .A1(ipA3[26]), .A2(n395), .Y(N222) );
  AND2X1_RVT U316 ( .A1(ipA3[25]), .A2(n393), .Y(N221) );
  AND2X1_RVT U317 ( .A1(ipA3[24]), .A2(n394), .Y(N220) );
  AND2X1_RVT U318 ( .A1(ipA1[18]), .A2(n395), .Y(N22) );
  AND2X1_RVT U319 ( .A1(ipA3[23]), .A2(n393), .Y(N219) );
  AND2X1_RVT U320 ( .A1(ipA3[22]), .A2(n394), .Y(N218) );
  AND2X1_RVT U321 ( .A1(ipA3[21]), .A2(n395), .Y(N217) );
  AND2X1_RVT U322 ( .A1(ipA3[20]), .A2(n393), .Y(N216) );
  AND2X1_RVT U323 ( .A1(ipA3[19]), .A2(n394), .Y(N215) );
  AND2X1_RVT U324 ( .A1(ipA3[18]), .A2(n395), .Y(N214) );
  AND2X1_RVT U325 ( .A1(ipA3[17]), .A2(n393), .Y(N213) );
  AND2X1_RVT U326 ( .A1(ipA3[16]), .A2(n394), .Y(N212) );
  AND2X1_RVT U327 ( .A1(ipA3[15]), .A2(n395), .Y(N211) );
  AND2X1_RVT U328 ( .A1(ipA3[14]), .A2(n393), .Y(N210) );
  AND2X1_RVT U329 ( .A1(ipA1[17]), .A2(n394), .Y(N21) );
  AND2X1_RVT U330 ( .A1(ipA3[13]), .A2(n395), .Y(N209) );
  AND2X1_RVT U331 ( .A1(ipA3[12]), .A2(n393), .Y(N208) );
  AND2X1_RVT U332 ( .A1(ipA3[11]), .A2(n394), .Y(N207) );
  AND2X1_RVT U333 ( .A1(ipA3[10]), .A2(n395), .Y(N206) );
  AND2X1_RVT U334 ( .A1(ipA3[9]), .A2(n394), .Y(N205) );
  AND2X1_RVT U335 ( .A1(ipA3[8]), .A2(n395), .Y(N204) );
  AND2X1_RVT U336 ( .A1(ipA3[7]), .A2(n393), .Y(N203) );
  AND2X1_RVT U337 ( .A1(ipA3[6]), .A2(n394), .Y(N202) );
  AND2X1_RVT U338 ( .A1(ipA3[5]), .A2(n395), .Y(N201) );
  AND2X1_RVT U339 ( .A1(ipA3[4]), .A2(n393), .Y(N200) );
  AND2X1_RVT U340 ( .A1(ipA1[16]), .A2(n394), .Y(N20) );
  AND2X1_RVT U341 ( .A1(ipA3[3]), .A2(n395), .Y(N199) );
  AND2X1_RVT U342 ( .A1(ipA3[2]), .A2(n393), .Y(N198) );
  AND2X1_RVT U343 ( .A1(ipA3[1]), .A2(n394), .Y(N197) );
  AND2X1_RVT U344 ( .A1(ipA3[0]), .A2(n395), .Y(N196) );
  AND2X1_RVT U345 ( .A1(ipA1[15]), .A2(n393), .Y(N19) );
  AND2X1_RVT U346 ( .A1(ipA1[14]), .A2(n394), .Y(N18) );
  AND2X1_RVT U347 ( .A1(ipA1[13]), .A2(n395), .Y(N17) );
  AND2X1_RVT U348 ( .A1(ipB2[31]), .A2(n393), .Y(N163) );
  AND2X1_RVT U349 ( .A1(ipB2[30]), .A2(n394), .Y(N162) );
  AND2X1_RVT U350 ( .A1(ipB2[29]), .A2(n395), .Y(N161) );
  AND2X1_RVT U351 ( .A1(ipB2[28]), .A2(n393), .Y(N160) );
  AND2X1_RVT U352 ( .A1(ipA1[12]), .A2(n394), .Y(N16) );
  AND2X1_RVT U353 ( .A1(ipB2[27]), .A2(n395), .Y(N159) );
  AND2X1_RVT U354 ( .A1(ipB2[26]), .A2(n391), .Y(N158) );
  AND2X1_RVT U355 ( .A1(ipB2[25]), .A2(n392), .Y(N157) );
  AND2X1_RVT U356 ( .A1(ipB2[24]), .A2(n395), .Y(N156) );
  AND2X1_RVT U357 ( .A1(ipB2[23]), .A2(n391), .Y(N155) );
  AND2X1_RVT U358 ( .A1(ipB2[22]), .A2(n392), .Y(N154) );
  AND2X1_RVT U359 ( .A1(ipB2[21]), .A2(n413), .Y(N153) );
  AND2X1_RVT U360 ( .A1(ipB2[20]), .A2(n391), .Y(N152) );
  AND2X1_RVT U361 ( .A1(ipB2[19]), .A2(n392), .Y(N151) );
  AND2X1_RVT U362 ( .A1(ipB2[18]), .A2(n414), .Y(N150) );
  AND2X1_RVT U363 ( .A1(ipA1[11]), .A2(n391), .Y(N15) );
  AND2X1_RVT U364 ( .A1(ipB2[17]), .A2(n392), .Y(N149) );
  AND2X1_RVT U365 ( .A1(ipB2[16]), .A2(n415), .Y(N148) );
  AND2X1_RVT U366 ( .A1(ipB2[15]), .A2(n391), .Y(N147) );
  AND2X1_RVT U367 ( .A1(ipB2[14]), .A2(n392), .Y(N146) );
  AND2X1_RVT U368 ( .A1(ipB2[13]), .A2(n411), .Y(N145) );
  AND2X1_RVT U369 ( .A1(ipB2[12]), .A2(n391), .Y(N144) );
  AND2X1_RVT U370 ( .A1(ipB2[11]), .A2(n392), .Y(N143) );
  AND2X1_RVT U371 ( .A1(ipB2[10]), .A2(n415), .Y(N142) );
  AND2X1_RVT U372 ( .A1(ipB2[9]), .A2(n391), .Y(N141) );
  AND2X1_RVT U373 ( .A1(ipB2[8]), .A2(n392), .Y(N140) );
  AND2X1_RVT U374 ( .A1(ipA1[10]), .A2(n411), .Y(N14) );
  AND2X1_RVT U375 ( .A1(ipB2[7]), .A2(n391), .Y(N139) );
  AND2X1_RVT U376 ( .A1(ipB2[6]), .A2(n392), .Y(N138) );
  AND2X1_RVT U377 ( .A1(ipB2[5]), .A2(n413), .Y(N137) );
  AND2X1_RVT U378 ( .A1(ipB2[4]), .A2(n391), .Y(N136) );
  AND2X1_RVT U379 ( .A1(ipB2[3]), .A2(n392), .Y(N135) );
  AND2X1_RVT U380 ( .A1(ipB2[2]), .A2(n414), .Y(N134) );
  AND2X1_RVT U381 ( .A1(ipB2[1]), .A2(n391), .Y(N133) );
  AND2X1_RVT U382 ( .A1(ipB2[0]), .A2(n392), .Y(N132) );
  AND2X1_RVT U383 ( .A1(ipA1[9]), .A2(n411), .Y(N13) );
  AND2X1_RVT U384 ( .A1(ipA1[8]), .A2(n391), .Y(N12) );
  AND2X1_RVT U385 ( .A1(ipA1[7]), .A2(n392), .Y(N11) );
  AND2X1_RVT U386 ( .A1(ipA1[6]), .A2(n393), .Y(N10) );
  OSPE_0 ospe00 ( .clk(clk), .rstnPipe(n409), .rstnPsum(rstnPsum[0]), .ipA(
        ipA0), .ipB(ipB0), .opA(opA00), .opB(opB00), .opC(opC00) );
  OSPE_15 ospe01 ( .clk(clk), .rstnPipe(n408), .rstnPsum(rstnPsum[1]), .ipA(
        opA00), .ipB(ipB1_d1), .opA(opA01), .opB(opB01), .opC(opC01) );
  OSPE_14 ospe02 ( .clk(clk), .rstnPipe(n385), .rstnPsum(rstnPsum[2]), .ipA(
        opA01), .ipB(ipB2_d2), .opA(opA02), .opB(opB02), .opC(opC02) );
  OSPE_13 ospe03 ( .clk(clk), .rstnPipe(n385), .rstnPsum(rstnPsum[3]), .ipA(
        opA02), .ipB(ipB3_d3), .opA({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32}), .opB(opB03), .opC(opC03) );
  OSPE_12 ospe10 ( .clk(clk), .rstnPipe(n385), .rstnPsum(rstnPsum[4]), .ipA(
        ipA1_d1), .ipB(opB00), .opA(opA10), .opB(opB10), .opC(opC10) );
  OSPE_11 ospe11 ( .clk(clk), .rstnPipe(n385), .rstnPsum(rstnPsum[5]), .ipA(
        opA10), .ipB(opB01), .opA(opA11), .opB(opB11), .opC(opC11) );
  OSPE_10 ospe12 ( .clk(clk), .rstnPipe(n408), .rstnPsum(rstnPsum[6]), .ipA(
        opA11), .ipB(opB02), .opA(opA12), .opB(opB12), .opC(opC12) );
  OSPE_9 ospe13 ( .clk(clk), .rstnPipe(n410), .rstnPsum(rstnPsum[7]), .ipA(
        opA12), .ipB(opB03), .opA({SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64}), .opB(opB13), .opC(opC13) );
  OSPE_8 ospe20 ( .clk(clk), .rstnPipe(n409), .rstnPsum(rstnPsum[8]), .ipA(
        ipA2_d2), .ipB(opB10), .opA(opA20), .opB(opB20), .opC(opC20) );
  OSPE_7 ospe21 ( .clk(clk), .rstnPipe(n408), .rstnPsum(rstnPsum[9]), .ipA(
        opA20), .ipB(opB11), .opA(opA21), .opB(opB21), .opC(opC21) );
  OSPE_6 ospe22 ( .clk(clk), .rstnPipe(n409), .rstnPsum(rstnPsum[10]), .ipA(
        opA21), .ipB(opB12), .opA(opA22), .opB(opB22), .opC(opC22) );
  OSPE_5 ospe23 ( .clk(clk), .rstnPipe(n410), .rstnPsum(rstnPsum[11]), .ipA(
        opA22), .ipB(opB13), .opA({SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96}), .opB(opB23), .opC(opC23) );
  OSPE_4 ospe30 ( .clk(clk), .rstnPipe(n409), .rstnPsum(rstnPsum[12]), .ipA(
        ipA3_d3), .ipB(opB20), .opA(opA30), .opB({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128}), .opC(opC30) );
  OSPE_3 ospe31 ( .clk(clk), .rstnPipe(n413), .rstnPsum(rstnPsum[13]), .ipA(
        opA30), .ipB(opB21), .opA(opA31), .opB({SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160}), .opC(opC31) );
  OSPE_2 ospe32 ( .clk(clk), .rstnPipe(n414), .rstnPsum(rstnPsum[14]), .ipA(
        opA31), .ipB(opB22), .opA(opA32), .opB({SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192}), .opC(opC32) );
  OSPE_1 ospe33 ( .clk(clk), .rstnPipe(n415), .rstnPsum(rstnPsum[15]), .ipA(
        opA32), .ipB(opB23), .opA({SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224}), .opB({SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256}), .opC(opC33) );
  DFFX1_RVT ipA1_d1_reg_31_ ( .D(N35), .CLK(clk), .Q(ipA1_d1[31]) );
  DFFX1_RVT ipA1_d1_reg_30_ ( .D(N34), .CLK(clk), .Q(ipA1_d1[30]) );
  DFFX1_RVT ipA1_d1_reg_29_ ( .D(N33), .CLK(clk), .Q(ipA1_d1[29]) );
  DFFX1_RVT ipA1_d1_reg_21_ ( .D(N25), .CLK(clk), .Q(ipA1_d1[21]) );
  DFFX1_RVT ipA1_d1_reg_28_ ( .D(N32), .CLK(clk), .Q(ipA1_d1[28]) );
  DFFX1_RVT ipA1_d1_reg_27_ ( .D(N31), .CLK(clk), .Q(ipA1_d1[27]) );
  DFFX1_RVT ipA1_d1_reg_26_ ( .D(N30), .CLK(clk), .Q(ipA1_d1[26]) );
  DFFX1_RVT ipA1_d1_reg_25_ ( .D(N29), .CLK(clk), .Q(ipA1_d1[25]) );
  DFFX1_RVT ipA1_d1_reg_24_ ( .D(N28), .CLK(clk), .Q(ipA1_d1[24]) );
  DFFX1_RVT ipA1_d1_reg_23_ ( .D(N27), .CLK(clk), .Q(ipA1_d1[23]) );
  DFFX1_RVT ipA1_d1_reg_22_ ( .D(N26), .CLK(clk), .Q(ipA1_d1[22]) );
  DFFX1_RVT ipA1_d1_reg_20_ ( .D(N24), .CLK(clk), .Q(ipA1_d1[20]) );
  DFFX1_RVT ipA1_d1_reg_19_ ( .D(N23), .CLK(clk), .Q(ipA1_d1[19]) );
  DFFX1_RVT ipA1_d1_reg_18_ ( .D(N22), .CLK(clk), .Q(ipA1_d1[18]) );
  DFFX1_RVT ipA1_d1_reg_17_ ( .D(N21), .CLK(clk), .Q(ipA1_d1[17]) );
  DFFX1_RVT ipA1_d1_reg_16_ ( .D(N20), .CLK(clk), .Q(ipA1_d1[16]) );
  DFFX1_RVT ipA1_d1_reg_15_ ( .D(N19), .CLK(clk), .Q(ipA1_d1[15]) );
  DFFX1_RVT ipA1_d1_reg_14_ ( .D(N18), .CLK(clk), .Q(ipA1_d1[14]) );
  DFFX1_RVT ipA1_d1_reg_13_ ( .D(N17), .CLK(clk), .Q(ipA1_d1[13]) );
  DFFX1_RVT ipA1_d1_reg_12_ ( .D(N16), .CLK(clk), .Q(ipA1_d1[12]) );
  DFFX1_RVT ipA1_d1_reg_11_ ( .D(N15), .CLK(clk), .Q(ipA1_d1[11]) );
  DFFX1_RVT ipA1_d1_reg_10_ ( .D(N14), .CLK(clk), .Q(ipA1_d1[10]) );
  DFFX1_RVT ipB1_d1_reg_15_ ( .D(N51), .CLK(clk), .Q(ipB1_d1[15]) );
  DFFX1_RVT ipB1_d1_reg_14_ ( .D(N50), .CLK(clk), .Q(ipB1_d1[14]) );
  DFFX1_RVT ipB1_d1_reg_13_ ( .D(N49), .CLK(clk), .Q(ipB1_d1[13]) );
  DFFX1_RVT ipB1_d1_reg_12_ ( .D(N48), .CLK(clk), .Q(ipB1_d1[12]) );
  DFFX1_RVT ipB1_d1_reg_11_ ( .D(N47), .CLK(clk), .Q(ipB1_d1[11]) );
  DFFX1_RVT ipB1_d1_reg_10_ ( .D(N46), .CLK(clk), .Q(ipB1_d1[10]) );
  DFFX1_RVT ipA1_d1_reg_9_ ( .D(N13), .CLK(clk), .Q(ipA1_d1[9]) );
  DFFX1_RVT ipA1_d1_reg_8_ ( .D(N12), .CLK(clk), .Q(ipA1_d1[8]) );
  DFFX1_RVT ipB1_d1_reg_9_ ( .D(N45), .CLK(clk), .Q(ipB1_d1[9]) );
  DFFX1_RVT ipB1_d1_reg_8_ ( .D(N44), .CLK(clk), .Q(ipB1_d1[8]) );
  DFFX1_RVT ipB1_d1_reg_7_ ( .D(N43), .CLK(clk), .Q(ipB1_d1[7]) );
  DFFX1_RVT ipB1_d1_reg_6_ ( .D(N42), .CLK(clk), .Q(ipB1_d1[6]) );
  DFFX1_RVT ipB1_d1_reg_5_ ( .D(N41), .CLK(clk), .Q(ipB1_d1[5]) );
  DFFX1_RVT ipA1_d1_reg_7_ ( .D(N11), .CLK(clk), .Q(ipA1_d1[7]) );
  DFFX1_RVT ipA1_d1_reg_6_ ( .D(N10), .CLK(clk), .Q(ipA1_d1[6]) );
  DFFX1_RVT ipA1_d1_reg_5_ ( .D(N9), .CLK(clk), .Q(ipA1_d1[5]) );
  DFFX1_RVT ipA1_d1_reg_4_ ( .D(N8), .CLK(clk), .Q(ipA1_d1[4]) );
  DFFX1_RVT ipB1_d1_reg_2_ ( .D(N38), .CLK(clk), .Q(ipB1_d1[2]) );
  DFFX1_RVT ipB1_d1_reg_1_ ( .D(N37), .CLK(clk), .Q(ipB1_d1[1]) );
  DFFX1_RVT ipB1_d1_reg_0_ ( .D(N36), .CLK(clk), .Q(ipB1_d1[0]) );
  DFFX1_RVT ipB1_d1_reg_31_ ( .D(N67), .CLK(clk), .Q(ipB1_d1[31]) );
  DFFX1_RVT ipB1_d1_reg_20_ ( .D(N56), .CLK(clk), .Q(ipB1_d1[20]) );
  DFFX1_RVT ipB1_d1_reg_19_ ( .D(N55), .CLK(clk), .Q(ipB1_d1[19]) );
  DFFX1_RVT ipB1_d1_reg_30_ ( .D(N66), .CLK(clk), .Q(ipB1_d1[30]) );
  DFFX1_RVT ipB1_d1_reg_18_ ( .D(N54), .CLK(clk), .Q(ipB1_d1[18]) );
  DFFX1_RVT ipB1_d1_reg_17_ ( .D(N53), .CLK(clk), .Q(ipB1_d1[17]) );
  DFFX1_RVT ipB1_d1_reg_16_ ( .D(N52), .CLK(clk), .Q(ipB1_d1[16]) );
  DFFX1_RVT ipB1_d1_reg_29_ ( .D(N65), .CLK(clk), .Q(ipB1_d1[29]) );
  DFFX1_RVT ipA1_d1_reg_3_ ( .D(N7), .CLK(clk), .Q(ipA1_d1[3]) );
  DFFX1_RVT ipA1_d1_reg_2_ ( .D(N6), .CLK(clk), .Q(ipA1_d1[2]) );
  DFFX1_RVT ipA1_d1_reg_1_ ( .D(N5), .CLK(clk), .Q(ipA1_d1[1]) );
  DFFX1_RVT ipA1_d1_reg_0_ ( .D(N4), .CLK(clk), .Q(ipA1_d1[0]) );
  DFFX1_RVT ipB1_d1_reg_4_ ( .D(N40), .CLK(clk), .Q(ipB1_d1[4]) );
  DFFX1_RVT ipB1_d1_reg_3_ ( .D(N39), .CLK(clk), .Q(ipB1_d1[3]) );
  DFFX1_RVT ipB1_d1_reg_28_ ( .D(N64), .CLK(clk), .Q(ipB1_d1[28]) );
  DFFX1_RVT ipB1_d1_reg_27_ ( .D(N63), .CLK(clk), .Q(ipB1_d1[27]) );
  DFFX1_RVT ipB1_d1_reg_26_ ( .D(N62), .CLK(clk), .Q(ipB1_d1[26]) );
  DFFX1_RVT ipB1_d1_reg_25_ ( .D(N61), .CLK(clk), .Q(ipB1_d1[25]) );
  DFFX1_RVT ipB1_d1_reg_24_ ( .D(N60), .CLK(clk), .Q(ipB1_d1[24]) );
  DFFX1_RVT ipB1_d1_reg_23_ ( .D(N59), .CLK(clk), .Q(ipB1_d1[23]) );
  DFFX1_RVT ipB1_d1_reg_22_ ( .D(N58), .CLK(clk), .Q(ipB1_d1[22]) );
  DFFX1_RVT ipB1_d1_reg_21_ ( .D(N57), .CLK(clk), .Q(ipB1_d1[21]) );
  DFFX1_RVT ipA2_d1_reg_31_ ( .D(N99), .CLK(clk), .QN(n384) );
  DFFX1_RVT ipA2_d1_reg_30_ ( .D(N98), .CLK(clk), .QN(n383) );
  DFFX1_RVT ipA2_d1_reg_29_ ( .D(N97), .CLK(clk), .QN(n382) );
  DFFX1_RVT ipA2_d1_reg_28_ ( .D(N96), .CLK(clk), .QN(n381) );
  DFFX1_RVT ipA2_d1_reg_27_ ( .D(N95), .CLK(clk), .QN(n380) );
  DFFX1_RVT ipA2_d1_reg_26_ ( .D(N94), .CLK(clk), .QN(n379) );
  DFFX1_RVT ipA2_d1_reg_25_ ( .D(N93), .CLK(clk), .QN(n378) );
  DFFX1_RVT ipA2_d1_reg_24_ ( .D(N92), .CLK(clk), .QN(n377) );
  DFFX1_RVT ipA2_d1_reg_23_ ( .D(N91), .CLK(clk), .QN(n376) );
  DFFX1_RVT ipA2_d1_reg_22_ ( .D(N90), .CLK(clk), .QN(n375) );
  DFFX1_RVT ipA2_d1_reg_21_ ( .D(N89), .CLK(clk), .QN(n374) );
  DFFX1_RVT ipA2_d1_reg_20_ ( .D(N88), .CLK(clk), .QN(n373) );
  DFFX1_RVT ipA2_d1_reg_19_ ( .D(N87), .CLK(clk), .QN(n372) );
  DFFX1_RVT ipA2_d1_reg_18_ ( .D(N86), .CLK(clk), .QN(n371) );
  DFFX1_RVT ipA2_d1_reg_17_ ( .D(N85), .CLK(clk), .QN(n370) );
  DFFX1_RVT ipA2_d1_reg_16_ ( .D(N84), .CLK(clk), .QN(n369) );
  DFFX1_RVT ipA2_d1_reg_15_ ( .D(N83), .CLK(clk), .QN(n368) );
  DFFX1_RVT ipA2_d1_reg_14_ ( .D(N82), .CLK(clk), .QN(n367) );
  DFFX1_RVT ipA2_d1_reg_13_ ( .D(N81), .CLK(clk), .QN(n366) );
  DFFX1_RVT ipA2_d1_reg_12_ ( .D(N80), .CLK(clk), .QN(n365) );
  DFFX1_RVT ipA2_d1_reg_11_ ( .D(N79), .CLK(clk), .QN(n364) );
  DFFX1_RVT ipA2_d1_reg_10_ ( .D(N78), .CLK(clk), .QN(n363) );
  DFFX1_RVT ipA2_d1_reg_9_ ( .D(N77), .CLK(clk), .QN(n362) );
  DFFX1_RVT ipA2_d1_reg_8_ ( .D(N76), .CLK(clk), .QN(n361) );
  DFFX1_RVT ipA2_d1_reg_7_ ( .D(N75), .CLK(clk), .QN(n360) );
  DFFX1_RVT ipA2_d1_reg_6_ ( .D(N74), .CLK(clk), .QN(n359) );
  DFFX1_RVT ipA2_d1_reg_5_ ( .D(N73), .CLK(clk), .QN(n358) );
  DFFX1_RVT ipA2_d1_reg_4_ ( .D(N72), .CLK(clk), .QN(n357) );
  DFFX1_RVT ipA2_d1_reg_3_ ( .D(N71), .CLK(clk), .QN(n356) );
  DFFX1_RVT ipA2_d1_reg_2_ ( .D(N70), .CLK(clk), .QN(n355) );
  DFFX1_RVT ipA2_d1_reg_1_ ( .D(N69), .CLK(clk), .QN(n354) );
  DFFX1_RVT ipA2_d1_reg_0_ ( .D(N68), .CLK(clk), .QN(n353) );
  DFFX1_RVT ipB2_d1_reg_31_ ( .D(N163), .CLK(clk), .QN(n320) );
  DFFX1_RVT ipB2_d1_reg_30_ ( .D(N162), .CLK(clk), .QN(n319) );
  DFFX1_RVT ipB2_d1_reg_29_ ( .D(N161), .CLK(clk), .QN(n318) );
  DFFX1_RVT ipB2_d1_reg_28_ ( .D(N160), .CLK(clk), .QN(n317) );
  DFFX1_RVT ipB2_d1_reg_27_ ( .D(N159), .CLK(clk), .QN(n316) );
  DFFX1_RVT ipB2_d1_reg_26_ ( .D(N158), .CLK(clk), .QN(n315) );
  DFFX1_RVT ipB2_d1_reg_25_ ( .D(N157), .CLK(clk), .QN(n314) );
  DFFX1_RVT ipB2_d1_reg_24_ ( .D(N156), .CLK(clk), .QN(n313) );
  DFFX1_RVT ipB2_d1_reg_23_ ( .D(N155), .CLK(clk), .QN(n312) );
  DFFX1_RVT ipB2_d1_reg_22_ ( .D(N154), .CLK(clk), .QN(n311) );
  DFFX1_RVT ipB2_d1_reg_21_ ( .D(N153), .CLK(clk), .QN(n310) );
  DFFX1_RVT ipB2_d1_reg_20_ ( .D(N152), .CLK(clk), .QN(n309) );
  DFFX1_RVT ipB2_d1_reg_19_ ( .D(N151), .CLK(clk), .QN(n308) );
  DFFX1_RVT ipB2_d1_reg_18_ ( .D(N150), .CLK(clk), .QN(n307) );
  DFFX1_RVT ipB2_d1_reg_17_ ( .D(N149), .CLK(clk), .QN(n306) );
  DFFX1_RVT ipB2_d1_reg_16_ ( .D(N148), .CLK(clk), .QN(n305) );
  DFFX1_RVT ipB2_d1_reg_15_ ( .D(N147), .CLK(clk), .QN(n304) );
  DFFX1_RVT ipB2_d1_reg_14_ ( .D(N146), .CLK(clk), .QN(n303) );
  DFFX1_RVT ipB2_d1_reg_13_ ( .D(N145), .CLK(clk), .QN(n302) );
  DFFX1_RVT ipB2_d1_reg_12_ ( .D(N144), .CLK(clk), .QN(n301) );
  DFFX1_RVT ipB2_d1_reg_11_ ( .D(N143), .CLK(clk), .QN(n300) );
  DFFX1_RVT ipB2_d1_reg_10_ ( .D(N142), .CLK(clk), .QN(n299) );
  DFFX1_RVT ipB2_d1_reg_9_ ( .D(N141), .CLK(clk), .QN(n298) );
  DFFX1_RVT ipB2_d1_reg_8_ ( .D(N140), .CLK(clk), .QN(n297) );
  DFFX1_RVT ipB2_d1_reg_7_ ( .D(N139), .CLK(clk), .QN(n296) );
  DFFX1_RVT ipB2_d1_reg_6_ ( .D(N138), .CLK(clk), .QN(n295) );
  DFFX1_RVT ipB2_d1_reg_5_ ( .D(N137), .CLK(clk), .QN(n294) );
  DFFX1_RVT ipB2_d1_reg_4_ ( .D(N136), .CLK(clk), .QN(n293) );
  DFFX1_RVT ipB2_d1_reg_3_ ( .D(N135), .CLK(clk), .QN(n292) );
  DFFX1_RVT ipB2_d1_reg_2_ ( .D(N134), .CLK(clk), .QN(n291) );
  DFFX1_RVT ipB2_d1_reg_1_ ( .D(N133), .CLK(clk), .QN(n290) );
  DFFX1_RVT ipB2_d1_reg_0_ ( .D(N132), .CLK(clk), .QN(n289) );
  DFFX1_RVT ipA3_d1_reg_31_ ( .D(N227), .CLK(clk), .QN(n256) );
  DFFX1_RVT ipA3_d1_reg_30_ ( .D(N226), .CLK(clk), .QN(n255) );
  DFFX1_RVT ipA3_d1_reg_29_ ( .D(N225), .CLK(clk), .QN(n254) );
  DFFX1_RVT ipA3_d1_reg_28_ ( .D(N224), .CLK(clk), .QN(n253) );
  DFFX1_RVT ipA3_d1_reg_27_ ( .D(N223), .CLK(clk), .QN(n252) );
  DFFX1_RVT ipA3_d1_reg_26_ ( .D(N222), .CLK(clk), .QN(n251) );
  DFFX1_RVT ipA3_d1_reg_25_ ( .D(N221), .CLK(clk), .QN(n250) );
  DFFX1_RVT ipA3_d1_reg_24_ ( .D(N220), .CLK(clk), .QN(n249) );
  DFFX1_RVT ipA3_d1_reg_23_ ( .D(N219), .CLK(clk), .QN(n248) );
  DFFX1_RVT ipA3_d1_reg_22_ ( .D(N218), .CLK(clk), .QN(n247) );
  DFFX1_RVT ipA3_d1_reg_21_ ( .D(N217), .CLK(clk), .QN(n246) );
  DFFX1_RVT ipA3_d1_reg_20_ ( .D(N216), .CLK(clk), .QN(n245) );
  DFFX1_RVT ipA3_d1_reg_19_ ( .D(N215), .CLK(clk), .QN(n244) );
  DFFX1_RVT ipA3_d1_reg_18_ ( .D(N214), .CLK(clk), .QN(n243) );
  DFFX1_RVT ipA3_d1_reg_17_ ( .D(N213), .CLK(clk), .QN(n242) );
  DFFX1_RVT ipA3_d1_reg_16_ ( .D(N212), .CLK(clk), .QN(n241) );
  DFFX1_RVT ipA3_d1_reg_15_ ( .D(N211), .CLK(clk), .QN(n240) );
  DFFX1_RVT ipA3_d1_reg_14_ ( .D(N210), .CLK(clk), .QN(n239) );
  DFFX1_RVT ipA3_d1_reg_13_ ( .D(N209), .CLK(clk), .QN(n238) );
  DFFX1_RVT ipA3_d1_reg_12_ ( .D(N208), .CLK(clk), .QN(n237) );
  DFFX1_RVT ipA3_d1_reg_11_ ( .D(N207), .CLK(clk), .QN(n236) );
  DFFX1_RVT ipA3_d1_reg_10_ ( .D(N206), .CLK(clk), .QN(n235) );
  DFFX1_RVT ipA3_d1_reg_9_ ( .D(N205), .CLK(clk), .QN(n234) );
  DFFX1_RVT ipA3_d1_reg_8_ ( .D(N204), .CLK(clk), .QN(n233) );
  DFFX1_RVT ipA3_d1_reg_7_ ( .D(N203), .CLK(clk), .QN(n232) );
  DFFX1_RVT ipA3_d1_reg_6_ ( .D(N202), .CLK(clk), .QN(n231) );
  DFFX1_RVT ipA3_d1_reg_5_ ( .D(N201), .CLK(clk), .QN(n230) );
  DFFX1_RVT ipA3_d1_reg_4_ ( .D(N200), .CLK(clk), .QN(n229) );
  DFFX1_RVT ipA3_d1_reg_3_ ( .D(N199), .CLK(clk), .QN(n228) );
  DFFX1_RVT ipA3_d1_reg_2_ ( .D(N198), .CLK(clk), .QN(n227) );
  DFFX1_RVT ipA3_d1_reg_1_ ( .D(N197), .CLK(clk), .QN(n226) );
  DFFX1_RVT ipA3_d1_reg_0_ ( .D(N196), .CLK(clk), .QN(n225) );
  DFFX1_RVT ipB3_d1_reg_31_ ( .D(N323), .CLK(clk), .QN(n128) );
  DFFX1_RVT ipB3_d1_reg_30_ ( .D(N322), .CLK(clk), .QN(n124) );
  DFFX1_RVT ipB3_d1_reg_29_ ( .D(N321), .CLK(clk), .QN(n120) );
  DFFX1_RVT ipB3_d1_reg_28_ ( .D(N320), .CLK(clk), .QN(n116) );
  DFFX1_RVT ipB3_d1_reg_27_ ( .D(N319), .CLK(clk), .QN(n112) );
  DFFX1_RVT ipB3_d1_reg_26_ ( .D(N318), .CLK(clk), .QN(n108) );
  DFFX1_RVT ipB3_d1_reg_25_ ( .D(N317), .CLK(clk), .QN(n104) );
  DFFX1_RVT ipB3_d1_reg_24_ ( .D(N316), .CLK(clk), .QN(n100) );
  DFFX1_RVT ipB3_d1_reg_23_ ( .D(N315), .CLK(clk), .QN(n96) );
  DFFX1_RVT ipB3_d1_reg_22_ ( .D(N314), .CLK(clk), .QN(n92) );
  DFFX1_RVT ipB3_d1_reg_21_ ( .D(N313), .CLK(clk), .QN(n88) );
  DFFX1_RVT ipB3_d1_reg_20_ ( .D(N312), .CLK(clk), .QN(n84) );
  DFFX1_RVT ipB3_d1_reg_19_ ( .D(N311), .CLK(clk), .QN(n80) );
  DFFX1_RVT ipB3_d1_reg_18_ ( .D(N310), .CLK(clk), .QN(n76) );
  DFFX1_RVT ipB3_d1_reg_17_ ( .D(N309), .CLK(clk), .QN(n72) );
  DFFX1_RVT ipB3_d1_reg_16_ ( .D(N308), .CLK(clk), .QN(n68) );
  DFFX1_RVT ipB3_d1_reg_15_ ( .D(N307), .CLK(clk), .QN(n64) );
  DFFX1_RVT ipB3_d1_reg_14_ ( .D(N306), .CLK(clk), .QN(n60) );
  DFFX1_RVT ipB3_d1_reg_13_ ( .D(N305), .CLK(clk), .QN(n56) );
  DFFX1_RVT ipB3_d1_reg_12_ ( .D(N304), .CLK(clk), .QN(n52) );
  DFFX1_RVT ipB3_d1_reg_11_ ( .D(N303), .CLK(clk), .QN(n48) );
  DFFX1_RVT ipB3_d1_reg_10_ ( .D(N302), .CLK(clk), .QN(n44) );
  DFFX1_RVT ipB3_d1_reg_9_ ( .D(N301), .CLK(clk), .QN(n40) );
  DFFX1_RVT ipB3_d1_reg_8_ ( .D(N300), .CLK(clk), .QN(n36) );
  DFFX1_RVT ipB3_d1_reg_7_ ( .D(N299), .CLK(clk), .QN(n32) );
  DFFX1_RVT ipB3_d1_reg_6_ ( .D(N298), .CLK(clk), .QN(n28) );
  DFFX1_RVT ipB3_d1_reg_5_ ( .D(N297), .CLK(clk), .QN(n24) );
  DFFX1_RVT ipB3_d1_reg_4_ ( .D(N296), .CLK(clk), .QN(n20) );
  DFFX1_RVT ipB3_d1_reg_3_ ( .D(N295), .CLK(clk), .QN(n16) );
  DFFX1_RVT ipB3_d1_reg_2_ ( .D(N294), .CLK(clk), .QN(n12) );
  DFFX1_RVT ipB3_d1_reg_1_ ( .D(N293), .CLK(clk), .QN(n8) );
  DFFX1_RVT ipB3_d1_reg_0_ ( .D(N292), .CLK(clk), .QN(n4) );
  INVX0_RVT U387 ( .A(n416), .Y(n409) );
  INVX0_RVT U388 ( .A(n416), .Y(n413) );
  INVX0_RVT U389 ( .A(n416), .Y(n414) );
  INVX0_RVT U390 ( .A(rstnPipe), .Y(n416) );
  INVX0_RVT U391 ( .A(n416), .Y(n408) );
  INVX1_RVT U392 ( .A(n416), .Y(n410) );
  INVX1_RVT U393 ( .A(n416), .Y(n411) );
  INVX1_RVT U394 ( .A(n416), .Y(n415) );
  INVX1_RVT U395 ( .A(n416), .Y(n412) );
  NBUFFX2_RVT U396 ( .A(n412), .Y(n385) );
  NBUFFX2_RVT U397 ( .A(n411), .Y(n386) );
  NBUFFX2_RVT U398 ( .A(n412), .Y(n387) );
  NBUFFX2_RVT U399 ( .A(n412), .Y(n388) );
  NBUFFX2_RVT U400 ( .A(rstnPipe), .Y(n389) );
  NBUFFX2_RVT U401 ( .A(n411), .Y(n390) );
  NBUFFX2_RVT U402 ( .A(n411), .Y(n391) );
  NBUFFX2_RVT U403 ( .A(n411), .Y(n392) );
  NBUFFX2_RVT U404 ( .A(n411), .Y(n393) );
  NBUFFX2_RVT U405 ( .A(n411), .Y(n394) );
  NBUFFX2_RVT U406 ( .A(n412), .Y(n395) );
  NBUFFX2_RVT U407 ( .A(n412), .Y(n396) );
  NBUFFX2_RVT U408 ( .A(n412), .Y(n397) );
  NBUFFX2_RVT U409 ( .A(n412), .Y(n398) );
  NBUFFX2_RVT U410 ( .A(n413), .Y(n399) );
  NBUFFX2_RVT U411 ( .A(n413), .Y(n400) );
  NBUFFX2_RVT U412 ( .A(n413), .Y(n401) );
  NBUFFX2_RVT U413 ( .A(n414), .Y(n402) );
  NBUFFX2_RVT U414 ( .A(n414), .Y(n403) );
  NBUFFX2_RVT U415 ( .A(n414), .Y(n404) );
  NBUFFX2_RVT U416 ( .A(n415), .Y(n405) );
  NBUFFX2_RVT U417 ( .A(n415), .Y(n406) );
  NBUFFX2_RVT U418 ( .A(n415), .Y(n407) );
endmodule


module DATA_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1_RVT U1 ( .A1(carry[9]), .A2(A[9]), .Y(SUM[9]) );
  INVX0_RVT U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DATA ( clk, rstnPipe, rstnAddr, addrInc, rstnPsum, latCnt, MemOutputA0, 
        MemOutputA1, MemOutputA2, MemOutputA3, MemOutputB0, MemOutputB1, 
        MemOutputB2, MemOutputB3, OpC00, OpC01, OpC02, OpC03, OpC10, OpC11, 
        OpC12, OpC13, OpC20, OpC21, OpC22, OpC23, OpC30, OpC31, OpC32, OpC33, 
        BankAddr );
  input [15:0] rstnPsum;
  input [3:0] latCnt;
  input [255:0] MemOutputA0;
  input [255:0] MemOutputA1;
  input [255:0] MemOutputA2;
  input [255:0] MemOutputA3;
  input [255:0] MemOutputB0;
  input [255:0] MemOutputB1;
  input [255:0] MemOutputB2;
  input [255:0] MemOutputB3;
  output [31:0] OpC00;
  output [31:0] OpC01;
  output [31:0] OpC02;
  output [31:0] OpC03;
  output [31:0] OpC10;
  output [31:0] OpC11;
  output [31:0] OpC12;
  output [31:0] OpC13;
  output [31:0] OpC20;
  output [31:0] OpC21;
  output [31:0] OpC22;
  output [31:0] OpC23;
  output [31:0] OpC30;
  output [31:0] OpC31;
  output [31:0] OpC32;
  output [31:0] OpC33;
  output [9:0] BankAddr;
  input clk, rstnPipe, rstnAddr, addrInc;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, opC11_d3_6_, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503,
         N504, N505, N506, N507, N508, N509, N510, N511, N512, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825,
         N826, N827, N828, N829, N830, N831, N832, N930, N931, N932, N933,
         N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944,
         N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955,
         N956, N957, N958, N959, N960, N999, N1057, N1058, N1059, N1060, N1061,
         N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071,
         N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081,
         N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1185, N1186, N1187,
         N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197,
         N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207,
         N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1281,
         N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291,
         N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301,
         N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311,
         N1312, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385,
         N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395,
         N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405,
         N1406, N1407, N1408, N1473, N1474, N1475, N1476, N1477, N1478, N1479,
         N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489,
         N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499,
         N1500, N1501, N1502, N1503, N1504, N1569, N1570, N1571, N1572, N1573,
         N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583,
         N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593,
         N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1633, N1634, N1635,
         N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645,
         N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655,
         N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1697,
         N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707,
         N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717,
         N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727,
         N1728, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769,
         N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779,
         N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789,
         N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799,
         N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, N1809,
         N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819,
         N1820, N1821, N1822, N1823, N1824, n2, n3, n6, n7, n8, n9, n10, n11,
         n13, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n401, n405, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n441, n445, n449, n453,
         n457, n461, n465, n469, n473, n477, n478, n479, n480, n481, n485,
         n489, n493, n497, n501, n505, n509, n513, n517, n521, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n929, n933, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1037, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1107, n1109, n1111, n1113, n1115,
         n1117, n1119, n1121, n1123, n1125, n1127, n1129, n1131, n1133, n1135,
         n1137, n1139, n1141, n1143, n1145, n1147, n1149, n1151, n1153, n1155,
         n1157, n1159, n1161, n1163, n1165, n1167, n1169, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1331, n1333, n1335, n1337, n1339, n1341, n1343, n1345, n1347,
         n1349, n1351, n1353, n1355, n1357, n1359, n1361, n1363, n1365, n1367,
         n1369, n1371, n1373, n1375, n1377, n1379, n1381, n1383, n1385, n1387,
         n1389, n1391, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1459, n1461, n1463, n1465, n1467,
         n1469, n1471, n1473, n1475, n1477, n1479, n1481, n1483, n1485, n1487,
         n1489, n1491, n1493, n1495, n1497, n1499, n1501, n1503, n1505, n1507,
         n1509, n1511, n1513, n1515, n1517, n1519, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1587,
         n1589, n1591, n1593, n1595, n1597, n1599, n1601, n1603, n1605, n1607,
         n1609, n1611, n1613, n1615, n1617, n1619, n1621, n1623, n1625, n1627,
         n1629, n1631, n1633, n1635, n1637, n1639, n1641, n1643, n1645, n1647,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1715, n1717, n1719, n1721, n1723, n1725, n1727,
         n1729, n1731, n1733, n1735, n1737, n1739, n1741, n1743, n1745, n1747,
         n1749, n1751, n1753, n1755, n1757, n1759, n1761, n1763, n1765, n1767,
         n1769, n1771, n1773, n1775, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1843, n1845, n1847,
         n1849, n1851, n1853, n1855, n1857, n1859, n1861, n1863, n1865, n1867,
         n1869, n1871, n1873, n1875, n1877, n1879, n1881, n1883, n1885, n1887,
         n1889, n1891, n1893, n1895, n1897, n1899, n1901, n1903, n1905, n1907,
         n1909, n1911, n1913, n1915, n1917, n1919, n1921, n1923, n1925, n1927,
         n1929, n1931, n1933, n1935, n1937, n1939, n1941, n1943, n1945, n1947,
         n1949, n1951, n1953, n1955, n1957, n1959, n1961, n1963, n1965, n1967,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2035, n2037, n2039, n2041, n2043, n2045, n2046,
         n2048, n2050, n2052, n2054, n2056, n2058, n2060, n2062, n2064, n2066,
         n2068, n2070, n2072, n2074, n2076, n2078, n2080, n2082, n2084, n2086,
         n2088, n2090, n2092, n2094, n2096, n2098, n2100, n2102, n2104, n2106,
         n2108, n2111, n2113, n2115, n2117, n2119, n2121, n2123, n2125, n2127,
         n2129, n2131, n2133, n2135, n2137, n2139, n2141, n2143, n2145, n2147,
         n2149, n2151, n2153, n2155, n2157, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2225, n2227,
         n2229, n2231, n2233, n2235, n2237, n2239, n2241, n2243, n2245, n2247,
         n2249, n2251, n2253, n2255, n2257, n2259, n2261, n2263, n2265, n2267,
         n2269, n2271, n2273, n2275, n2277, n2279, n2281, n2283, n2285, n2287,
         n2289, n2291, n2293, n2295, n2297, n2299, n2301, n2303, n2305, n2307,
         n2309, n2311, n2313, n2315, n2317, n2319, n2321, n2323, n2325, n2327,
         n2329, n2331, n2333, n2335, n2337, n2339, n2341, n2343, n2345, n2347,
         n2349, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2417, n2419, n2421, n2423, n2425, n2427,
         n2429, n2431, n2433, n2435, n2437, n2439, n2441, n2443, n2445, n2447,
         n2449, n2451, n2453, n2455, n2457, n2459, n2461, n2463, n2465, n2467,
         n2469, n2471, n2473, n2475, n2477, n2479, n2481, n2483, n2485, n2487,
         n2489, n2491, n2493, n2495, n2497, n2499, n2501, n2503, n2505, n2507,
         n2509, n2511, n2513, n2515, n2517, n2519, n2521, n2523, n2525, n2527,
         n2529, n2531, n2533, n2535, n2537, n2539, n2541, n2543, n2545, n2547,
         n2549, n2551, n2553, n2555, n2557, n2559, n2561, n2563, n2565, n2567,
         n2569, n2571, n2573, n2575, n2577, n2579, n2581, n2583, n2585, n2587,
         n2589, n2591, n2593, n2595, n2597, n2599, n2601, n2603, n2605, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2673, n2675, n2677, n2679, n2681, n2683, n2685, n2687,
         n2689, n2691, n2693, n2695, n2697, n2699, n2701, n2703, n2705, n2707,
         n2709, n2711, n2713, n2715, n2717, n2719, n2721, n2723, n2725, n2727,
         n2729, n2731, n2733, n2735, n2737, n2739, n2741, n2743, n2745, n2747,
         n2749, n2751, n2753, n2755, n2757, n2759, n2761, n2763, n2765, n2767,
         n2769, n2771, n2773, n2775, n2777, n2779, n2781, n2783, n2785, n2787,
         n2789, n2791, n2793, n2795, n2797, n2799, n2801, n2803, n2805, n2807,
         n2809, n2811, n2813, n2815, n2817, n2819, n2821, n2823, n2825, n2827,
         n2829, n2831, n2833, n2835, n2837, n2839, n2841, n2843, n2845, n2847,
         n2849, n2851, n2853, n2855, n2857, n2859, n2861, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2929, n2931, n2933, n2935, n2937, n2939, n2941, n2943, n2945, n2947,
         n2949, n2951, n2953, n2955, n2957, n2959, n2961, n2963, n2965, n2967,
         n2969, n2971, n2973, n2975, n2977, n2979, n2981, n2983, n2985, n2987,
         n2989, n2991, n2993, n2995, n2997, n2999, n3001, n3003, n3005, n3007,
         n3009, n3011, n3013, n3015, n3017, n3019, n3021, n3023, n3025, n3027,
         n3029, n3031, n3033, n3035, n3037, n3039, n3041, n3043, n3045, n3047,
         n3049, n3051, n3053, n3055, n3057, n3059, n3061, n3063, n3065, n3067,
         n3069, n3071, n3073, n3075, n3077, n3079, n3081, n3083, n3085, n3087,
         n3089, n3091, n3093, n3095, n3097, n3099, n3101, n3103, n3105, n3107,
         n3109, n3111, n3113, n3115, n3117, n3119, n3121, n3123, n3125, n3127,
         n3129, n3131, n3133, n3135, n3137, n3139, n3141, n3143, n3145, n3147,
         n3149, n3151, n3153, n3155, n3157, n3159, n3161, n3163, n3165, n3167,
         n3169, n3171, n3173, n3175, n3177, n3179, n3181, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n1, n4, n5, n12, n14, n15, n16, n398, n399, n400, n402, n403, n404,
         n406, n407, n408, n418, n419, n420, n438, n439, n440, n442, n443,
         n444, n450, n451, n452, n454, n455, n456, n458, n459, n460, n462,
         n463, n464, n466, n467, n468, n470, n471, n472, n474, n475, n476,
         n482, n483, n484, n486, n487, n488, n490, n491, n492, n494, n495,
         n496, n498, n499, n500, n502, n503, n504, n506, n507, n508, n510,
         n511, n512, n514, n515, n516, n518, n519, n520, n522, n523, n524,
         n926, n927, n928, n930, n931, n932, n934, n935, n936, n946, n947,
         n948, n990, n991, n992, n1034, n1035, n1036, n1038, n1039, n1040,
         n1041, n1112, n3180, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574;
  wire   [31:0] ipA0;
  wire   [31:0] ipA1;
  wire   [31:0] ipA2;
  wire   [31:0] ipA3;
  wire   [31:0] ipB0;
  wire   [31:0] ipB1;
  wire   [31:0] ipB2;
  wire   [31:0] ipB3;
  wire   [31:0] opC00_out;
  wire   [31:0] opC01_out;
  wire   [31:0] opC02_out;
  wire   [31:0] opC03_out;
  wire   [31:0] opC10_out;
  wire   [31:0] opC11_out;
  wire   [31:0] opC12_out;
  wire   [31:0] opC13_out;
  wire   [31:0] opC20_out;
  wire   [31:0] opC21_out;
  wire   [31:0] opC22_out;
  wire   [31:0] opC23_out;
  wire   [31:0] opC30_out;
  wire   [31:0] opC31_out;
  wire   [31:0] opC32_out;

  SDFFX1_RVT opC00_d5_reg_31_ ( .D(n3449), .SI(1'b0), .SE(n1074), .CLK(clk), 
        .QN(n3183) );
  SDFFX1_RVT opC00_d5_reg_29_ ( .D(n3441), .SI(1'b0), .SE(n1076), .CLK(clk), 
        .QN(n3179) );
  SDFFX1_RVT opC00_d5_reg_28_ ( .D(n3441), .SI(1'b0), .SE(n1077), .CLK(clk), 
        .QN(n3177) );
  SDFFX1_RVT opC00_d5_reg_27_ ( .D(n3441), .SI(1'b0), .SE(n1078), .CLK(clk), 
        .QN(n3175) );
  SDFFX1_RVT opC00_d5_reg_26_ ( .D(n3459), .SI(1'b0), .SE(n1079), .CLK(clk), 
        .QN(n3173) );
  SDFFX1_RVT opC00_d5_reg_25_ ( .D(n3460), .SI(1'b0), .SE(n1080), .CLK(clk), 
        .QN(n3171) );
  SDFFX1_RVT opC00_d5_reg_24_ ( .D(n3464), .SI(1'b0), .SE(n1081), .CLK(clk), 
        .QN(n3169) );
  SDFFX1_RVT opC00_d5_reg_23_ ( .D(n3465), .SI(1'b0), .SE(n1082), .CLK(clk), 
        .QN(n3167) );
  SDFFX1_RVT opC00_d5_reg_22_ ( .D(n3442), .SI(1'b0), .SE(n1083), .CLK(clk), 
        .QN(n3165) );
  SDFFX1_RVT opC00_d5_reg_21_ ( .D(n3478), .SI(1'b0), .SE(n1084), .CLK(clk), 
        .QN(n3163) );
  SDFFX1_RVT opC00_d5_reg_20_ ( .D(n3446), .SI(1'b0), .SE(n1085), .CLK(clk), 
        .QN(n3161) );
  SDFFX1_RVT opC00_d5_reg_19_ ( .D(n3447), .SI(1'b0), .SE(n1086), .CLK(clk), 
        .QN(n3159) );
  SDFFX1_RVT opC00_d5_reg_18_ ( .D(n3451), .SI(1'b0), .SE(n1087), .CLK(clk), 
        .QN(n3157) );
  SDFFX1_RVT opC00_d5_reg_17_ ( .D(n3452), .SI(1'b0), .SE(n1088), .CLK(clk), 
        .QN(n3155) );
  SDFFX1_RVT opC00_d5_reg_16_ ( .D(n3461), .SI(1'b0), .SE(n1089), .CLK(clk), 
        .QN(n3153) );
  SDFFX1_RVT opC00_d5_reg_15_ ( .D(n3448), .SI(1'b0), .SE(n1090), .CLK(clk), 
        .QN(n3151) );
  SDFFX1_RVT opC00_d5_reg_14_ ( .D(n3450), .SI(1'b0), .SE(n1091), .CLK(clk), 
        .QN(n3149) );
  SDFFX1_RVT opC00_d5_reg_13_ ( .D(n3442), .SI(1'b0), .SE(n1092), .CLK(clk), 
        .QN(n3147) );
  SDFFX1_RVT opC00_d5_reg_12_ ( .D(n3445), .SI(1'b0), .SE(n1093), .CLK(clk), 
        .QN(n3145) );
  SDFFX1_RVT opC00_d5_reg_11_ ( .D(n3472), .SI(1'b0), .SE(n1094), .CLK(clk), 
        .QN(n3143) );
  SDFFX1_RVT opC00_d5_reg_10_ ( .D(n3474), .SI(1'b0), .SE(n1095), .CLK(clk), 
        .QN(n3141) );
  SDFFX1_RVT opC00_d5_reg_9_ ( .D(n3462), .SI(1'b0), .SE(n1096), .CLK(clk), 
        .QN(n3139) );
  SDFFX1_RVT opC00_d5_reg_8_ ( .D(n3461), .SI(1'b0), .SE(n1097), .CLK(clk), 
        .QN(n3137) );
  SDFFX1_RVT opC00_d5_reg_7_ ( .D(n3463), .SI(1'b0), .SE(n1098), .CLK(clk), 
        .QN(n3135) );
  SDFFX1_RVT opC00_d5_reg_6_ ( .D(n3456), .SI(1'b0), .SE(n1099), .CLK(clk), 
        .QN(n3133) );
  SDFFX1_RVT opC00_d5_reg_5_ ( .D(n3458), .SI(1'b0), .SE(n1100), .CLK(clk), 
        .QN(n3131) );
  SDFFX1_RVT opC00_d5_reg_4_ ( .D(n3442), .SI(1'b0), .SE(n1101), .CLK(clk), 
        .QN(n3129) );
  SDFFX1_RVT opC00_d5_reg_3_ ( .D(n3477), .SI(1'b0), .SE(n1102), .CLK(clk), 
        .QN(n3127) );
  SDFFX1_RVT opC00_d5_reg_2_ ( .D(n3479), .SI(1'b0), .SE(n1103), .CLK(clk), 
        .QN(n3125) );
  SDFFX1_RVT opC00_d5_reg_1_ ( .D(n3480), .SI(1'b0), .SE(n1104), .CLK(clk), 
        .QN(n3123) );
  SDFFX1_RVT opC00_d5_reg_0_ ( .D(n3466), .SI(1'b0), .SE(n1105), .CLK(clk), 
        .QN(n3121) );
  SDFFX1_RVT opC00_d4_reg_31_ ( .D(n3481), .SI(1'b0), .SE(n3183), .CLK(clk), 
        .QN(n3119) );
  SDFFX1_RVT opC00_d4_reg_30_ ( .D(n3449), .SI(1'b0), .SE(n3181), .CLK(clk), 
        .QN(n3117) );
  SDFFX1_RVT opC00_d4_reg_29_ ( .D(n3458), .SI(1'b0), .SE(n3179), .CLK(clk), 
        .QN(n3115) );
  SDFFX1_RVT opC00_d4_reg_28_ ( .D(n3453), .SI(1'b0), .SE(n3177), .CLK(clk), 
        .QN(n3113) );
  SDFFX1_RVT opC00_d4_reg_27_ ( .D(n3454), .SI(1'b0), .SE(n3175), .CLK(clk), 
        .QN(n3111) );
  SDFFX1_RVT opC00_d4_reg_26_ ( .D(n3443), .SI(1'b0), .SE(n3173), .CLK(clk), 
        .QN(n3109) );
  SDFFX1_RVT opC00_d4_reg_25_ ( .D(n3476), .SI(1'b0), .SE(n3171), .CLK(clk), 
        .QN(n3107) );
  SDFFX1_RVT opC00_d4_reg_24_ ( .D(n3475), .SI(1'b0), .SE(n3169), .CLK(clk), 
        .QN(n3105) );
  SDFFX1_RVT opC00_d4_reg_23_ ( .D(n3457), .SI(1'b0), .SE(n3167), .CLK(clk), 
        .QN(n3103) );
  SDFFX1_RVT opC00_d4_reg_22_ ( .D(n3455), .SI(1'b0), .SE(n3165), .CLK(clk), 
        .QN(n3101) );
  SDFFX1_RVT opC00_d4_reg_21_ ( .D(n3464), .SI(1'b0), .SE(n3163), .CLK(clk), 
        .QN(n3099) );
  SDFFX1_RVT opC00_d4_reg_20_ ( .D(n3367), .SI(1'b0), .SE(n3161), .CLK(clk), 
        .QN(n3097) );
  SDFFX1_RVT opC00_d4_reg_19_ ( .D(n3454), .SI(1'b0), .SE(n3159), .CLK(clk), 
        .QN(n3095) );
  SDFFX1_RVT opC00_d4_reg_18_ ( .D(n3465), .SI(1'b0), .SE(n3157), .CLK(clk), 
        .QN(n3093) );
  SDFFX1_RVT opC00_d4_reg_17_ ( .D(n3443), .SI(1'b0), .SE(n3155), .CLK(clk), 
        .QN(n3091) );
  SDFFX1_RVT opC00_d4_reg_16_ ( .D(n3440), .SI(1'b0), .SE(n3153), .CLK(clk), 
        .QN(n3089) );
  SDFFX1_RVT opC00_d4_reg_15_ ( .D(n3440), .SI(1'b0), .SE(n3151), .CLK(clk), 
        .QN(n3087) );
  SDFFX1_RVT opC00_d4_reg_14_ ( .D(n3440), .SI(1'b0), .SE(n3149), .CLK(clk), 
        .QN(n3085) );
  SDFFX1_RVT opC00_d4_reg_13_ ( .D(n3440), .SI(1'b0), .SE(n3147), .CLK(clk), 
        .QN(n3083) );
  SDFFX1_RVT opC00_d4_reg_12_ ( .D(n3440), .SI(1'b0), .SE(n3145), .CLK(clk), 
        .QN(n3081) );
  SDFFX1_RVT opC00_d4_reg_11_ ( .D(n3440), .SI(1'b0), .SE(n3143), .CLK(clk), 
        .QN(n3079) );
  SDFFX1_RVT opC00_d4_reg_10_ ( .D(n3440), .SI(1'b0), .SE(n3141), .CLK(clk), 
        .QN(n3077) );
  SDFFX1_RVT opC00_d4_reg_9_ ( .D(n3440), .SI(1'b0), .SE(n3139), .CLK(clk), 
        .QN(n3075) );
  SDFFX1_RVT opC00_d4_reg_8_ ( .D(n3440), .SI(1'b0), .SE(n3137), .CLK(clk), 
        .QN(n3073) );
  SDFFX1_RVT opC00_d4_reg_7_ ( .D(n3440), .SI(1'b0), .SE(n3135), .CLK(clk), 
        .QN(n3071) );
  SDFFX1_RVT opC00_d4_reg_6_ ( .D(n3440), .SI(1'b0), .SE(n3133), .CLK(clk), 
        .QN(n3069) );
  SDFFX1_RVT opC00_d4_reg_5_ ( .D(n3440), .SI(1'b0), .SE(n3131), .CLK(clk), 
        .QN(n3067) );
  SDFFX1_RVT opC00_d4_reg_4_ ( .D(n3440), .SI(1'b0), .SE(n3129), .CLK(clk), 
        .QN(n3065) );
  SDFFX1_RVT opC00_d4_reg_3_ ( .D(n3440), .SI(1'b0), .SE(n3127), .CLK(clk), 
        .QN(n3063) );
  SDFFX1_RVT opC00_d4_reg_2_ ( .D(n3439), .SI(1'b0), .SE(n3125), .CLK(clk), 
        .QN(n3061) );
  SDFFX1_RVT opC00_d4_reg_1_ ( .D(n3439), .SI(1'b0), .SE(n3123), .CLK(clk), 
        .QN(n3059) );
  SDFFX1_RVT opC00_d4_reg_0_ ( .D(n3439), .SI(1'b0), .SE(n3121), .CLK(clk), 
        .QN(n3057) );
  SDFFX1_RVT opC00_d3_reg_31_ ( .D(n3439), .SI(1'b0), .SE(n3119), .CLK(clk), 
        .QN(n3055) );
  SDFFX1_RVT opC00_d3_reg_30_ ( .D(n3439), .SI(1'b0), .SE(n3117), .CLK(clk), 
        .QN(n3053) );
  SDFFX1_RVT opC00_d3_reg_29_ ( .D(n3439), .SI(1'b0), .SE(n3115), .CLK(clk), 
        .QN(n3051) );
  SDFFX1_RVT opC00_d3_reg_28_ ( .D(n3439), .SI(1'b0), .SE(n3113), .CLK(clk), 
        .QN(n3049) );
  SDFFX1_RVT opC00_d3_reg_27_ ( .D(n3439), .SI(1'b0), .SE(n3111), .CLK(clk), 
        .QN(n3047) );
  SDFFX1_RVT opC00_d3_reg_26_ ( .D(n3439), .SI(1'b0), .SE(n3109), .CLK(clk), 
        .QN(n3045) );
  SDFFX1_RVT opC00_d3_reg_25_ ( .D(n3439), .SI(1'b0), .SE(n3107), .CLK(clk), 
        .QN(n3043) );
  SDFFX1_RVT opC00_d3_reg_24_ ( .D(n3439), .SI(1'b0), .SE(n3105), .CLK(clk), 
        .QN(n3041) );
  SDFFX1_RVT opC00_d3_reg_23_ ( .D(n3439), .SI(1'b0), .SE(n3103), .CLK(clk), 
        .QN(n3039) );
  SDFFX1_RVT opC00_d3_reg_22_ ( .D(n3473), .SI(1'b0), .SE(n3101), .CLK(clk), 
        .QN(n3037) );
  SDFFX1_RVT opC00_d3_reg_21_ ( .D(n3346), .SI(1'b0), .SE(n3099), .CLK(clk), 
        .QN(n3035) );
  SDFFX1_RVT opC00_d3_reg_20_ ( .D(n3370), .SI(1'b0), .SE(n3097), .CLK(clk), 
        .QN(n3033) );
  SDFFX1_RVT opC00_d3_reg_19_ ( .D(n3442), .SI(1'b0), .SE(n3095), .CLK(clk), 
        .QN(n3031) );
  SDFFX1_RVT opC00_d3_reg_18_ ( .D(n3478), .SI(1'b0), .SE(n3093), .CLK(clk), 
        .QN(n3029) );
  SDFFX1_RVT opC00_d3_reg_17_ ( .D(n3446), .SI(1'b0), .SE(n3091), .CLK(clk), 
        .QN(n3027) );
  SDFFX1_RVT opC00_d3_reg_16_ ( .D(n3447), .SI(1'b0), .SE(n3089), .CLK(clk), 
        .QN(n3025) );
  SDFFX1_RVT opC00_d3_reg_15_ ( .D(n3451), .SI(1'b0), .SE(n3087), .CLK(clk), 
        .QN(n3023) );
  SDFFX1_RVT opC00_d3_reg_14_ ( .D(n3452), .SI(1'b0), .SE(n3085), .CLK(clk), 
        .QN(n3021) );
  SDFFX1_RVT opC00_d3_reg_13_ ( .D(n3463), .SI(1'b0), .SE(n3083), .CLK(clk), 
        .QN(n3019) );
  SDFFX1_RVT opC00_d3_reg_12_ ( .D(n3448), .SI(1'b0), .SE(n3081), .CLK(clk), 
        .QN(n3017) );
  SDFFX1_RVT opC00_d3_reg_11_ ( .D(n3450), .SI(1'b0), .SE(n3079), .CLK(clk), 
        .QN(n3015) );
  SDFFX1_RVT opC00_d3_reg_10_ ( .D(n3444), .SI(1'b0), .SE(n3077), .CLK(clk), 
        .QN(n3013) );
  SDFFX1_RVT opC00_d3_reg_9_ ( .D(n3444), .SI(1'b0), .SE(n3075), .CLK(clk), 
        .QN(n3011) );
  SDFFX1_RVT opC00_d3_reg_8_ ( .D(n3438), .SI(1'b0), .SE(n3073), .CLK(clk), 
        .QN(n3009) );
  SDFFX1_RVT opC00_d3_reg_7_ ( .D(n3438), .SI(1'b0), .SE(n3071), .CLK(clk), 
        .QN(n3007) );
  SDFFX1_RVT opC00_d3_reg_6_ ( .D(n3438), .SI(1'b0), .SE(n3069), .CLK(clk), 
        .QN(n3005) );
  SDFFX1_RVT opC00_d3_reg_5_ ( .D(n3438), .SI(1'b0), .SE(n3067), .CLK(clk), 
        .QN(n3003) );
  SDFFX1_RVT opC00_d3_reg_4_ ( .D(n3438), .SI(1'b0), .SE(n3065), .CLK(clk), 
        .QN(n3001) );
  SDFFX1_RVT opC00_d3_reg_3_ ( .D(n3438), .SI(1'b0), .SE(n3063), .CLK(clk), 
        .QN(n2999) );
  SDFFX1_RVT opC00_d3_reg_2_ ( .D(n3438), .SI(1'b0), .SE(n3061), .CLK(clk), 
        .QN(n2997) );
  SDFFX1_RVT opC00_d3_reg_1_ ( .D(n3438), .SI(1'b0), .SE(n3059), .CLK(clk), 
        .QN(n2995) );
  SDFFX1_RVT opC00_d3_reg_0_ ( .D(n3438), .SI(1'b0), .SE(n3057), .CLK(clk), 
        .QN(n2993) );
  SDFFX1_RVT opC00_d2_reg_31_ ( .D(n3438), .SI(1'b0), .SE(n3055), .CLK(clk), 
        .QN(n2991) );
  SDFFX1_RVT opC00_d2_reg_30_ ( .D(n3438), .SI(1'b0), .SE(n3053), .CLK(clk), 
        .QN(n2989) );
  SDFFX1_RVT opC00_d2_reg_29_ ( .D(n3438), .SI(1'b0), .SE(n3051), .CLK(clk), 
        .QN(n2987) );
  SDFFX1_RVT opC00_d2_reg_28_ ( .D(n3438), .SI(1'b0), .SE(n3049), .CLK(clk), 
        .QN(n2985) );
  SDFFX1_RVT opC00_d2_reg_27_ ( .D(n3438), .SI(1'b0), .SE(n3047), .CLK(clk), 
        .QN(n2983) );
  SDFFX1_RVT opC00_d2_reg_26_ ( .D(n3437), .SI(1'b0), .SE(n3045), .CLK(clk), 
        .QN(n2981) );
  SDFFX1_RVT opC00_d2_reg_25_ ( .D(n3437), .SI(1'b0), .SE(n3043), .CLK(clk), 
        .QN(n2979) );
  SDFFX1_RVT opC00_d2_reg_24_ ( .D(n3437), .SI(1'b0), .SE(n3041), .CLK(clk), 
        .QN(n2977) );
  SDFFX1_RVT opC00_d2_reg_23_ ( .D(n3437), .SI(1'b0), .SE(n3039), .CLK(clk), 
        .QN(n2975) );
  SDFFX1_RVT opC00_d2_reg_22_ ( .D(n3437), .SI(1'b0), .SE(n3037), .CLK(clk), 
        .QN(n2973) );
  SDFFX1_RVT opC00_d2_reg_21_ ( .D(n3437), .SI(1'b0), .SE(n3035), .CLK(clk), 
        .QN(n2971) );
  SDFFX1_RVT opC00_d2_reg_20_ ( .D(n3437), .SI(1'b0), .SE(n3033), .CLK(clk), 
        .QN(n2969) );
  SDFFX1_RVT opC00_d2_reg_19_ ( .D(n3437), .SI(1'b0), .SE(n3031), .CLK(clk), 
        .QN(n2967) );
  SDFFX1_RVT opC00_d2_reg_18_ ( .D(n3437), .SI(1'b0), .SE(n3029), .CLK(clk), 
        .QN(n2965) );
  SDFFX1_RVT opC00_d2_reg_17_ ( .D(n3437), .SI(1'b0), .SE(n3027), .CLK(clk), 
        .QN(n2963) );
  SDFFX1_RVT opC00_d2_reg_16_ ( .D(n3437), .SI(1'b0), .SE(n3025), .CLK(clk), 
        .QN(n2961) );
  SDFFX1_RVT opC00_d2_reg_15_ ( .D(n3437), .SI(1'b0), .SE(n3023), .CLK(clk), 
        .QN(n2959) );
  SDFFX1_RVT opC00_d2_reg_14_ ( .D(n3437), .SI(1'b0), .SE(n3021), .CLK(clk), 
        .QN(n2957) );
  SDFFX1_RVT opC00_d2_reg_13_ ( .D(n3437), .SI(1'b0), .SE(n3019), .CLK(clk), 
        .QN(n2955) );
  SDFFX1_RVT opC00_d2_reg_12_ ( .D(n3436), .SI(1'b0), .SE(n3017), .CLK(clk), 
        .QN(n2953) );
  SDFFX1_RVT opC00_d2_reg_11_ ( .D(n3436), .SI(1'b0), .SE(n3015), .CLK(clk), 
        .QN(n2951) );
  SDFFX1_RVT opC00_d2_reg_10_ ( .D(n3436), .SI(1'b0), .SE(n3013), .CLK(clk), 
        .QN(n2949) );
  SDFFX1_RVT opC00_d2_reg_9_ ( .D(n3436), .SI(1'b0), .SE(n3011), .CLK(clk), 
        .QN(n2947) );
  SDFFX1_RVT opC00_d2_reg_8_ ( .D(n3436), .SI(1'b0), .SE(n3009), .CLK(clk), 
        .QN(n2945) );
  SDFFX1_RVT opC00_d2_reg_7_ ( .D(n3436), .SI(1'b0), .SE(n3007), .CLK(clk), 
        .QN(n2943) );
  SDFFX1_RVT opC00_d2_reg_6_ ( .D(n3436), .SI(1'b0), .SE(n3005), .CLK(clk), 
        .QN(n2941) );
  SDFFX1_RVT opC00_d2_reg_5_ ( .D(n3436), .SI(1'b0), .SE(n3003), .CLK(clk), 
        .QN(n2939) );
  SDFFX1_RVT opC00_d2_reg_4_ ( .D(n3436), .SI(1'b0), .SE(n3001), .CLK(clk), 
        .QN(n2937) );
  SDFFX1_RVT opC00_d2_reg_3_ ( .D(n3436), .SI(1'b0), .SE(n2999), .CLK(clk), 
        .QN(n2935) );
  SDFFX1_RVT opC00_d2_reg_2_ ( .D(n3436), .SI(1'b0), .SE(n2997), .CLK(clk), 
        .QN(n2933) );
  SDFFX1_RVT opC00_d2_reg_1_ ( .D(n3436), .SI(1'b0), .SE(n2995), .CLK(clk), 
        .QN(n2931) );
  SDFFX1_RVT opC00_d2_reg_0_ ( .D(n3436), .SI(1'b0), .SE(n2993), .CLK(clk), 
        .QN(n2929) );
  SDFFX1_RVT opC00_d1_reg_31_ ( .D(n3436), .SI(1'b0), .SE(n2991), .CLK(clk), 
        .Q(OpC00[31]) );
  SDFFX1_RVT opC00_d1_reg_30_ ( .D(n3460), .SI(1'b0), .SE(n2989), .CLK(clk), 
        .Q(OpC00[30]) );
  SDFFX1_RVT opC00_d1_reg_29_ ( .D(n3439), .SI(1'b0), .SE(n2987), .CLK(clk), 
        .Q(OpC00[29]) );
  SDFFX1_RVT opC00_d1_reg_28_ ( .D(n3418), .SI(1'b0), .SE(n2985), .CLK(clk), 
        .Q(OpC00[28]) );
  SDFFX1_RVT opC00_d1_reg_27_ ( .D(n3439), .SI(1'b0), .SE(n2983), .CLK(clk), 
        .Q(OpC00[27]) );
  SDFFX1_RVT opC00_d1_reg_26_ ( .D(n3453), .SI(1'b0), .SE(n2981), .CLK(clk), 
        .Q(OpC00[26]) );
  SDFFX1_RVT opC00_d1_reg_25_ ( .D(n3454), .SI(1'b0), .SE(n2979), .CLK(clk), 
        .Q(OpC00[25]) );
  SDFFX1_RVT opC00_d1_reg_24_ ( .D(n3445), .SI(1'b0), .SE(n2977), .CLK(clk), 
        .Q(OpC00[24]) );
  SDFFX1_RVT opC00_d1_reg_23_ ( .D(n3476), .SI(1'b0), .SE(n2975), .CLK(clk), 
        .Q(OpC00[23]) );
  SDFFX1_RVT opC00_d1_reg_22_ ( .D(n3475), .SI(1'b0), .SE(n2973), .CLK(clk), 
        .Q(OpC00[22]) );
  SDFFX1_RVT opC00_d1_reg_21_ ( .D(n3457), .SI(1'b0), .SE(n2971), .CLK(clk), 
        .Q(OpC00[21]) );
  SDFFX1_RVT opC00_d1_reg_20_ ( .D(n3455), .SI(1'b0), .SE(n2969), .CLK(clk), 
        .Q(OpC00[20]) );
  SDFFX1_RVT opC00_d1_reg_19_ ( .D(n3348), .SI(1'b0), .SE(n2967), .CLK(clk), 
        .Q(OpC00[19]) );
  SDFFX1_RVT opC00_d1_reg_18_ ( .D(n3367), .SI(1'b0), .SE(n2965), .CLK(clk), 
        .Q(OpC00[18]) );
  SDFFX1_RVT opC00_d1_reg_17_ ( .D(n3453), .SI(1'b0), .SE(n2963), .CLK(clk), 
        .Q(OpC00[17]) );
  SDFFX1_RVT opC00_d1_reg_16_ ( .D(n3465), .SI(1'b0), .SE(n2961), .CLK(clk), 
        .Q(OpC00[16]) );
  SDFFX1_RVT opC00_d1_reg_15_ ( .D(n3445), .SI(1'b0), .SE(n2959), .CLK(clk), 
        .Q(OpC00[15]) );
  SDFFX1_RVT opC00_d1_reg_14_ ( .D(n3435), .SI(1'b0), .SE(n2957), .CLK(clk), 
        .Q(OpC00[14]) );
  SDFFX1_RVT opC00_d1_reg_13_ ( .D(n3435), .SI(1'b0), .SE(n2955), .CLK(clk), 
        .Q(OpC00[13]) );
  SDFFX1_RVT opC00_d1_reg_12_ ( .D(n3435), .SI(1'b0), .SE(n2953), .CLK(clk), 
        .Q(OpC00[12]) );
  SDFFX1_RVT opC00_d1_reg_11_ ( .D(n3435), .SI(1'b0), .SE(n2951), .CLK(clk), 
        .Q(OpC00[11]) );
  SDFFX1_RVT opC00_d1_reg_10_ ( .D(n3435), .SI(1'b0), .SE(n2949), .CLK(clk), 
        .Q(OpC00[10]) );
  SDFFX1_RVT opC00_d1_reg_9_ ( .D(n3435), .SI(1'b0), .SE(n2947), .CLK(clk), 
        .Q(OpC00[9]) );
  SDFFX1_RVT opC00_d1_reg_8_ ( .D(n3435), .SI(1'b0), .SE(n2945), .CLK(clk), 
        .Q(OpC00[8]) );
  SDFFX1_RVT opC00_d1_reg_7_ ( .D(n3435), .SI(1'b0), .SE(n2943), .CLK(clk), 
        .Q(OpC00[7]) );
  SDFFX1_RVT opC00_d1_reg_6_ ( .D(n3435), .SI(1'b0), .SE(n2941), .CLK(clk), 
        .Q(OpC00[6]) );
  SDFFX1_RVT opC00_d1_reg_5_ ( .D(n3435), .SI(1'b0), .SE(n2939), .CLK(clk), 
        .Q(OpC00[5]) );
  SDFFX1_RVT opC00_d1_reg_4_ ( .D(n3435), .SI(1'b0), .SE(n2937), .CLK(clk), 
        .Q(OpC00[4]) );
  SDFFX1_RVT opC00_d1_reg_3_ ( .D(n3435), .SI(1'b0), .SE(n2935), .CLK(clk), 
        .Q(OpC00[3]) );
  SDFFX1_RVT opC00_d1_reg_2_ ( .D(n3435), .SI(1'b0), .SE(n2933), .CLK(clk), 
        .Q(OpC00[2]) );
  SDFFX1_RVT opC00_d1_reg_1_ ( .D(n3435), .SI(1'b0), .SE(n2931), .CLK(clk), 
        .Q(OpC00[1]) );
  SDFFX1_RVT opC00_d1_reg_0_ ( .D(n3434), .SI(1'b0), .SE(n2929), .CLK(clk), 
        .Q(OpC00[0]) );
  SDFFX1_RVT opC01_d4_reg_31_ ( .D(n3434), .SI(1'b0), .SE(n2895), .CLK(clk), 
        .QN(n2863) );
  SDFFX1_RVT opC01_d4_reg_30_ ( .D(n3434), .SI(1'b0), .SE(n2894), .CLK(clk), 
        .QN(n2861) );
  SDFFX1_RVT opC01_d4_reg_29_ ( .D(n3434), .SI(1'b0), .SE(n2893), .CLK(clk), 
        .QN(n2859) );
  SDFFX1_RVT opC01_d4_reg_28_ ( .D(n3434), .SI(1'b0), .SE(n2892), .CLK(clk), 
        .QN(n2857) );
  SDFFX1_RVT opC01_d4_reg_27_ ( .D(n3434), .SI(1'b0), .SE(n2891), .CLK(clk), 
        .QN(n2855) );
  SDFFX1_RVT opC01_d4_reg_26_ ( .D(n3434), .SI(1'b0), .SE(n2890), .CLK(clk), 
        .QN(n2853) );
  SDFFX1_RVT opC01_d4_reg_25_ ( .D(n3434), .SI(1'b0), .SE(n2889), .CLK(clk), 
        .QN(n2851) );
  SDFFX1_RVT opC01_d4_reg_24_ ( .D(n3434), .SI(1'b0), .SE(n2888), .CLK(clk), 
        .QN(n2849) );
  SDFFX1_RVT opC01_d4_reg_23_ ( .D(n3434), .SI(1'b0), .SE(n2887), .CLK(clk), 
        .QN(n2847) );
  SDFFX1_RVT opC01_d4_reg_22_ ( .D(n3434), .SI(1'b0), .SE(n2886), .CLK(clk), 
        .QN(n2845) );
  SDFFX1_RVT opC01_d4_reg_21_ ( .D(n3434), .SI(1'b0), .SE(n2885), .CLK(clk), 
        .QN(n2843) );
  SDFFX1_RVT opC01_d4_reg_20_ ( .D(n3434), .SI(1'b0), .SE(n2884), .CLK(clk), 
        .QN(n2841) );
  SDFFX1_RVT opC01_d4_reg_19_ ( .D(n3434), .SI(1'b0), .SE(n2883), .CLK(clk), 
        .QN(n2839) );
  SDFFX1_RVT opC01_d4_reg_18_ ( .D(n3433), .SI(1'b0), .SE(n2882), .CLK(clk), 
        .QN(n2837) );
  SDFFX1_RVT opC01_d4_reg_17_ ( .D(n3433), .SI(1'b0), .SE(n2881), .CLK(clk), 
        .QN(n2835) );
  SDFFX1_RVT opC01_d4_reg_16_ ( .D(n3433), .SI(1'b0), .SE(n2880), .CLK(clk), 
        .QN(n2833) );
  SDFFX1_RVT opC01_d4_reg_15_ ( .D(n3433), .SI(1'b0), .SE(n2879), .CLK(clk), 
        .QN(n2831) );
  SDFFX1_RVT opC01_d4_reg_14_ ( .D(n3433), .SI(1'b0), .SE(n2878), .CLK(clk), 
        .QN(n2829) );
  SDFFX1_RVT opC01_d4_reg_13_ ( .D(n3433), .SI(1'b0), .SE(n2877), .CLK(clk), 
        .QN(n2827) );
  SDFFX1_RVT opC01_d4_reg_12_ ( .D(n3433), .SI(1'b0), .SE(n2876), .CLK(clk), 
        .QN(n2825) );
  SDFFX1_RVT opC01_d4_reg_11_ ( .D(n3433), .SI(1'b0), .SE(n2875), .CLK(clk), 
        .QN(n2823) );
  SDFFX1_RVT opC01_d4_reg_10_ ( .D(n3433), .SI(1'b0), .SE(n2874), .CLK(clk), 
        .QN(n2821) );
  SDFFX1_RVT opC01_d4_reg_9_ ( .D(n3433), .SI(1'b0), .SE(n2873), .CLK(clk), 
        .QN(n2819) );
  SDFFX1_RVT opC01_d4_reg_8_ ( .D(n3433), .SI(1'b0), .SE(n2872), .CLK(clk), 
        .QN(n2817) );
  SDFFX1_RVT opC01_d4_reg_7_ ( .D(n3433), .SI(1'b0), .SE(n2871), .CLK(clk), 
        .QN(n2815) );
  SDFFX1_RVT opC01_d4_reg_6_ ( .D(n3433), .SI(1'b0), .SE(n2870), .CLK(clk), 
        .QN(n2813) );
  SDFFX1_RVT opC01_d4_reg_5_ ( .D(n3433), .SI(1'b0), .SE(n2869), .CLK(clk), 
        .QN(n2811) );
  SDFFX1_RVT opC01_d4_reg_4_ ( .D(n3432), .SI(1'b0), .SE(n2868), .CLK(clk), 
        .QN(n2809) );
  SDFFX1_RVT opC01_d4_reg_3_ ( .D(n3432), .SI(1'b0), .SE(n2867), .CLK(clk), 
        .QN(n2807) );
  SDFFX1_RVT opC01_d4_reg_2_ ( .D(n3432), .SI(1'b0), .SE(n2866), .CLK(clk), 
        .QN(n2805) );
  SDFFX1_RVT opC01_d4_reg_1_ ( .D(n3432), .SI(1'b0), .SE(n2865), .CLK(clk), 
        .QN(n2803) );
  SDFFX1_RVT opC01_d4_reg_0_ ( .D(n3432), .SI(1'b0), .SE(n2864), .CLK(clk), 
        .QN(n2801) );
  SDFFX1_RVT opC01_d3_reg_31_ ( .D(n3432), .SI(1'b0), .SE(n2863), .CLK(clk), 
        .QN(n2799) );
  SDFFX1_RVT opC01_d3_reg_30_ ( .D(n3432), .SI(1'b0), .SE(n2861), .CLK(clk), 
        .QN(n2797) );
  SDFFX1_RVT opC01_d3_reg_29_ ( .D(n3432), .SI(1'b0), .SE(n2859), .CLK(clk), 
        .QN(n2795) );
  SDFFX1_RVT opC01_d3_reg_28_ ( .D(n3432), .SI(1'b0), .SE(n2857), .CLK(clk), 
        .QN(n2793) );
  SDFFX1_RVT opC01_d3_reg_27_ ( .D(n3432), .SI(1'b0), .SE(n2855), .CLK(clk), 
        .QN(n2791) );
  SDFFX1_RVT opC01_d3_reg_26_ ( .D(n3432), .SI(1'b0), .SE(n2853), .CLK(clk), 
        .QN(n2789) );
  SDFFX1_RVT opC01_d3_reg_25_ ( .D(n3432), .SI(1'b0), .SE(n2851), .CLK(clk), 
        .QN(n2787) );
  SDFFX1_RVT opC01_d3_reg_24_ ( .D(n3431), .SI(1'b0), .SE(n2849), .CLK(clk), 
        .QN(n2785) );
  SDFFX1_RVT opC01_d3_reg_23_ ( .D(n3431), .SI(1'b0), .SE(n2847), .CLK(clk), 
        .QN(n2783) );
  SDFFX1_RVT opC01_d3_reg_22_ ( .D(n3431), .SI(1'b0), .SE(n2845), .CLK(clk), 
        .QN(n2781) );
  SDFFX1_RVT opC01_d3_reg_21_ ( .D(n3431), .SI(1'b0), .SE(n2843), .CLK(clk), 
        .QN(n2779) );
  SDFFX1_RVT opC01_d3_reg_20_ ( .D(n3431), .SI(1'b0), .SE(n2841), .CLK(clk), 
        .QN(n2777) );
  SDFFX1_RVT opC01_d3_reg_19_ ( .D(n3431), .SI(1'b0), .SE(n2839), .CLK(clk), 
        .QN(n2775) );
  SDFFX1_RVT opC01_d3_reg_18_ ( .D(n3431), .SI(1'b0), .SE(n2837), .CLK(clk), 
        .QN(n2773) );
  SDFFX1_RVT opC01_d3_reg_17_ ( .D(n3431), .SI(1'b0), .SE(n2835), .CLK(clk), 
        .QN(n2771) );
  SDFFX1_RVT opC01_d3_reg_16_ ( .D(n3431), .SI(1'b0), .SE(n2833), .CLK(clk), 
        .QN(n2769) );
  SDFFX1_RVT opC01_d3_reg_15_ ( .D(n3431), .SI(1'b0), .SE(n2831), .CLK(clk), 
        .QN(n2767) );
  SDFFX1_RVT opC01_d3_reg_14_ ( .D(n3431), .SI(1'b0), .SE(n2829), .CLK(clk), 
        .QN(n2765) );
  SDFFX1_RVT opC01_d3_reg_13_ ( .D(n3431), .SI(1'b0), .SE(n2827), .CLK(clk), 
        .QN(n2763) );
  SDFFX1_RVT opC01_d3_reg_12_ ( .D(n3431), .SI(1'b0), .SE(n2825), .CLK(clk), 
        .QN(n2761) );
  SDFFX1_RVT opC01_d3_reg_11_ ( .D(n3431), .SI(1'b0), .SE(n2823), .CLK(clk), 
        .QN(n2759) );
  SDFFX1_RVT opC01_d3_reg_10_ ( .D(n3430), .SI(1'b0), .SE(n2821), .CLK(clk), 
        .QN(n2757) );
  SDFFX1_RVT opC01_d3_reg_9_ ( .D(n3430), .SI(1'b0), .SE(n2819), .CLK(clk), 
        .QN(n2755) );
  SDFFX1_RVT opC01_d3_reg_8_ ( .D(n3430), .SI(1'b0), .SE(n2817), .CLK(clk), 
        .QN(n2753) );
  SDFFX1_RVT opC01_d3_reg_7_ ( .D(n3430), .SI(1'b0), .SE(n2815), .CLK(clk), 
        .QN(n2751) );
  SDFFX1_RVT opC01_d3_reg_6_ ( .D(n3430), .SI(1'b0), .SE(n2813), .CLK(clk), 
        .QN(n2749) );
  SDFFX1_RVT opC01_d3_reg_5_ ( .D(n3430), .SI(1'b0), .SE(n2811), .CLK(clk), 
        .QN(n2747) );
  SDFFX1_RVT opC01_d3_reg_4_ ( .D(n3430), .SI(1'b0), .SE(n2809), .CLK(clk), 
        .QN(n2745) );
  SDFFX1_RVT opC01_d3_reg_3_ ( .D(n3430), .SI(1'b0), .SE(n2807), .CLK(clk), 
        .QN(n2743) );
  SDFFX1_RVT opC01_d3_reg_2_ ( .D(n3430), .SI(1'b0), .SE(n2805), .CLK(clk), 
        .QN(n2741) );
  SDFFX1_RVT opC01_d3_reg_1_ ( .D(n3430), .SI(1'b0), .SE(n2803), .CLK(clk), 
        .QN(n2739) );
  SDFFX1_RVT opC01_d3_reg_0_ ( .D(n3430), .SI(1'b0), .SE(n2801), .CLK(clk), 
        .QN(n2737) );
  SDFFX1_RVT opC01_d2_reg_31_ ( .D(n3430), .SI(1'b0), .SE(n2799), .CLK(clk), 
        .QN(n2735) );
  SDFFX1_RVT opC01_d2_reg_30_ ( .D(n3430), .SI(1'b0), .SE(n2797), .CLK(clk), 
        .QN(n2733) );
  SDFFX1_RVT opC01_d2_reg_29_ ( .D(n3430), .SI(1'b0), .SE(n2795), .CLK(clk), 
        .QN(n2731) );
  SDFFX1_RVT opC01_d2_reg_28_ ( .D(n3429), .SI(1'b0), .SE(n2793), .CLK(clk), 
        .QN(n2729) );
  SDFFX1_RVT opC01_d2_reg_27_ ( .D(n3429), .SI(1'b0), .SE(n2791), .CLK(clk), 
        .QN(n2727) );
  SDFFX1_RVT opC01_d2_reg_26_ ( .D(n3429), .SI(1'b0), .SE(n2789), .CLK(clk), 
        .QN(n2725) );
  SDFFX1_RVT opC01_d2_reg_25_ ( .D(n3429), .SI(1'b0), .SE(n2787), .CLK(clk), 
        .QN(n2723) );
  SDFFX1_RVT opC01_d2_reg_24_ ( .D(n3429), .SI(1'b0), .SE(n2785), .CLK(clk), 
        .QN(n2721) );
  SDFFX1_RVT opC01_d2_reg_23_ ( .D(n3429), .SI(1'b0), .SE(n2783), .CLK(clk), 
        .QN(n2719) );
  SDFFX1_RVT opC01_d2_reg_22_ ( .D(n3429), .SI(1'b0), .SE(n2781), .CLK(clk), 
        .QN(n2717) );
  SDFFX1_RVT opC01_d2_reg_21_ ( .D(n3429), .SI(1'b0), .SE(n2779), .CLK(clk), 
        .QN(n2715) );
  SDFFX1_RVT opC01_d2_reg_20_ ( .D(n3429), .SI(1'b0), .SE(n2777), .CLK(clk), 
        .QN(n2713) );
  SDFFX1_RVT opC01_d2_reg_19_ ( .D(n3429), .SI(1'b0), .SE(n2775), .CLK(clk), 
        .QN(n2711) );
  SDFFX1_RVT opC01_d2_reg_18_ ( .D(n3429), .SI(1'b0), .SE(n2773), .CLK(clk), 
        .QN(n2709) );
  SDFFX1_RVT opC01_d2_reg_17_ ( .D(n3429), .SI(1'b0), .SE(n2771), .CLK(clk), 
        .QN(n2707) );
  SDFFX1_RVT opC01_d2_reg_16_ ( .D(n3429), .SI(1'b0), .SE(n2769), .CLK(clk), 
        .QN(n2705) );
  SDFFX1_RVT opC01_d2_reg_15_ ( .D(n3429), .SI(1'b0), .SE(n2767), .CLK(clk), 
        .QN(n2703) );
  SDFFX1_RVT opC01_d2_reg_14_ ( .D(n3428), .SI(1'b0), .SE(n2765), .CLK(clk), 
        .QN(n2701) );
  SDFFX1_RVT opC01_d2_reg_13_ ( .D(n3428), .SI(1'b0), .SE(n2763), .CLK(clk), 
        .QN(n2699) );
  SDFFX1_RVT opC01_d2_reg_12_ ( .D(n3428), .SI(1'b0), .SE(n2761), .CLK(clk), 
        .QN(n2697) );
  SDFFX1_RVT opC01_d2_reg_11_ ( .D(n3428), .SI(1'b0), .SE(n2759), .CLK(clk), 
        .QN(n2695) );
  SDFFX1_RVT opC01_d2_reg_10_ ( .D(n3428), .SI(1'b0), .SE(n2757), .CLK(clk), 
        .QN(n2693) );
  SDFFX1_RVT opC01_d2_reg_9_ ( .D(n3428), .SI(1'b0), .SE(n2755), .CLK(clk), 
        .QN(n2691) );
  SDFFX1_RVT opC01_d2_reg_8_ ( .D(n3428), .SI(1'b0), .SE(n2753), .CLK(clk), 
        .QN(n2689) );
  SDFFX1_RVT opC01_d2_reg_7_ ( .D(n3428), .SI(1'b0), .SE(n2751), .CLK(clk), 
        .QN(n2687) );
  SDFFX1_RVT opC01_d2_reg_6_ ( .D(n3428), .SI(1'b0), .SE(n2749), .CLK(clk), 
        .QN(n2685) );
  SDFFX1_RVT opC01_d2_reg_5_ ( .D(n3428), .SI(1'b0), .SE(n2747), .CLK(clk), 
        .QN(n2683) );
  SDFFX1_RVT opC01_d2_reg_4_ ( .D(n3428), .SI(1'b0), .SE(n2745), .CLK(clk), 
        .QN(n2681) );
  SDFFX1_RVT opC01_d2_reg_3_ ( .D(n3428), .SI(1'b0), .SE(n2743), .CLK(clk), 
        .QN(n2679) );
  SDFFX1_RVT opC01_d2_reg_2_ ( .D(n3428), .SI(1'b0), .SE(n2741), .CLK(clk), 
        .QN(n2677) );
  SDFFX1_RVT opC01_d2_reg_1_ ( .D(n3428), .SI(1'b0), .SE(n2739), .CLK(clk), 
        .QN(n2675) );
  SDFFX1_RVT opC01_d2_reg_0_ ( .D(n3427), .SI(1'b0), .SE(n2737), .CLK(clk), 
        .QN(n2673) );
  SDFFX1_RVT opC01_d1_reg_31_ ( .D(n3427), .SI(1'b0), .SE(n2735), .CLK(clk), 
        .Q(OpC01[31]) );
  SDFFX1_RVT opC01_d1_reg_30_ ( .D(n3427), .SI(1'b0), .SE(n2733), .CLK(clk), 
        .Q(OpC01[30]) );
  SDFFX1_RVT opC01_d1_reg_29_ ( .D(n3427), .SI(1'b0), .SE(n2731), .CLK(clk), 
        .Q(OpC01[29]) );
  SDFFX1_RVT opC01_d1_reg_28_ ( .D(n3427), .SI(1'b0), .SE(n2729), .CLK(clk), 
        .Q(OpC01[28]) );
  SDFFX1_RVT opC01_d1_reg_27_ ( .D(n3427), .SI(1'b0), .SE(n2727), .CLK(clk), 
        .Q(OpC01[27]) );
  SDFFX1_RVT opC01_d1_reg_26_ ( .D(n3427), .SI(1'b0), .SE(n2725), .CLK(clk), 
        .Q(OpC01[26]) );
  SDFFX1_RVT opC01_d1_reg_25_ ( .D(n3432), .SI(1'b0), .SE(n2723), .CLK(clk), 
        .Q(OpC01[25]) );
  SDFFX1_RVT opC01_d1_reg_24_ ( .D(n3432), .SI(1'b0), .SE(n2721), .CLK(clk), 
        .Q(OpC01[24]) );
  SDFFX1_RVT opC01_d1_reg_23_ ( .D(n3422), .SI(1'b0), .SE(n2719), .CLK(clk), 
        .Q(OpC01[23]) );
  SDFFX1_RVT opC01_d1_reg_22_ ( .D(n3427), .SI(1'b0), .SE(n2717), .CLK(clk), 
        .Q(OpC01[22]) );
  SDFFX1_RVT opC01_d1_reg_21_ ( .D(n3427), .SI(1'b0), .SE(n2715), .CLK(clk), 
        .Q(OpC01[21]) );
  SDFFX1_RVT opC01_d1_reg_20_ ( .D(n3427), .SI(1'b0), .SE(n2713), .CLK(clk), 
        .Q(OpC01[20]) );
  SDFFX1_RVT opC01_d1_reg_19_ ( .D(n3427), .SI(1'b0), .SE(n2711), .CLK(clk), 
        .Q(OpC01[19]) );
  SDFFX1_RVT opC01_d1_reg_18_ ( .D(n3426), .SI(1'b0), .SE(n2709), .CLK(clk), 
        .Q(OpC01[18]) );
  SDFFX1_RVT opC01_d1_reg_17_ ( .D(n3426), .SI(1'b0), .SE(n2707), .CLK(clk), 
        .Q(OpC01[17]) );
  SDFFX1_RVT opC01_d1_reg_16_ ( .D(n3426), .SI(1'b0), .SE(n2705), .CLK(clk), 
        .Q(OpC01[16]) );
  SDFFX1_RVT opC01_d1_reg_15_ ( .D(n3426), .SI(1'b0), .SE(n2703), .CLK(clk), 
        .Q(OpC01[15]) );
  SDFFX1_RVT opC01_d1_reg_14_ ( .D(n3426), .SI(1'b0), .SE(n2701), .CLK(clk), 
        .Q(OpC01[14]) );
  SDFFX1_RVT opC01_d1_reg_13_ ( .D(n3426), .SI(1'b0), .SE(n2699), .CLK(clk), 
        .Q(OpC01[13]) );
  SDFFX1_RVT opC01_d1_reg_12_ ( .D(n3426), .SI(1'b0), .SE(n2697), .CLK(clk), 
        .Q(OpC01[12]) );
  SDFFX1_RVT opC01_d1_reg_11_ ( .D(n3426), .SI(1'b0), .SE(n2695), .CLK(clk), 
        .Q(OpC01[11]) );
  SDFFX1_RVT opC01_d1_reg_10_ ( .D(n3426), .SI(1'b0), .SE(n2693), .CLK(clk), 
        .Q(OpC01[10]) );
  SDFFX1_RVT opC01_d1_reg_9_ ( .D(n3426), .SI(1'b0), .SE(n2691), .CLK(clk), 
        .Q(OpC01[9]) );
  SDFFX1_RVT opC01_d1_reg_8_ ( .D(n3426), .SI(1'b0), .SE(n2689), .CLK(clk), 
        .Q(OpC01[8]) );
  SDFFX1_RVT opC01_d1_reg_7_ ( .D(n3426), .SI(1'b0), .SE(n2687), .CLK(clk), 
        .Q(OpC01[7]) );
  SDFFX1_RVT opC01_d1_reg_6_ ( .D(n3426), .SI(1'b0), .SE(n2685), .CLK(clk), 
        .Q(OpC01[6]) );
  SDFFX1_RVT opC01_d1_reg_5_ ( .D(n3426), .SI(1'b0), .SE(n2683), .CLK(clk), 
        .Q(OpC01[5]) );
  SDFFX1_RVT opC01_d1_reg_4_ ( .D(n3425), .SI(1'b0), .SE(n2681), .CLK(clk), 
        .Q(OpC01[4]) );
  SDFFX1_RVT opC01_d1_reg_3_ ( .D(n3425), .SI(1'b0), .SE(n2679), .CLK(clk), 
        .Q(OpC01[3]) );
  SDFFX1_RVT opC01_d1_reg_2_ ( .D(n3425), .SI(1'b0), .SE(n2677), .CLK(clk), 
        .Q(OpC01[2]) );
  SDFFX1_RVT opC01_d1_reg_1_ ( .D(n3425), .SI(1'b0), .SE(n2675), .CLK(clk), 
        .Q(OpC01[1]) );
  SDFFX1_RVT opC01_d1_reg_0_ ( .D(n3425), .SI(1'b0), .SE(n2673), .CLK(clk), 
        .Q(OpC01[0]) );
  SDFFX1_RVT opC10_d4_reg_31_ ( .D(n3425), .SI(1'b0), .SE(n2639), .CLK(clk), 
        .QN(n2607) );
  SDFFX1_RVT opC10_d4_reg_30_ ( .D(n3425), .SI(1'b0), .SE(n2638), .CLK(clk), 
        .QN(n2605) );
  SDFFX1_RVT opC10_d4_reg_29_ ( .D(n3425), .SI(1'b0), .SE(n2637), .CLK(clk), 
        .QN(n2603) );
  SDFFX1_RVT opC10_d4_reg_28_ ( .D(n3425), .SI(1'b0), .SE(n2636), .CLK(clk), 
        .QN(n2601) );
  SDFFX1_RVT opC10_d4_reg_27_ ( .D(n3425), .SI(1'b0), .SE(n2635), .CLK(clk), 
        .QN(n2599) );
  SDFFX1_RVT opC10_d4_reg_26_ ( .D(n3425), .SI(1'b0), .SE(n2634), .CLK(clk), 
        .QN(n2597) );
  SDFFX1_RVT opC10_d4_reg_25_ ( .D(n3425), .SI(1'b0), .SE(n2633), .CLK(clk), 
        .QN(n2595) );
  SDFFX1_RVT opC10_d4_reg_24_ ( .D(n3425), .SI(1'b0), .SE(n2632), .CLK(clk), 
        .QN(n2593) );
  SDFFX1_RVT opC10_d4_reg_23_ ( .D(n3425), .SI(1'b0), .SE(n2631), .CLK(clk), 
        .QN(n2591) );
  SDFFX1_RVT opC10_d4_reg_22_ ( .D(n3424), .SI(1'b0), .SE(n2630), .CLK(clk), 
        .QN(n2589) );
  SDFFX1_RVT opC10_d4_reg_21_ ( .D(n3424), .SI(1'b0), .SE(n2629), .CLK(clk), 
        .QN(n2587) );
  SDFFX1_RVT opC10_d4_reg_20_ ( .D(n3424), .SI(1'b0), .SE(n2628), .CLK(clk), 
        .QN(n2585) );
  SDFFX1_RVT opC10_d4_reg_19_ ( .D(n3424), .SI(1'b0), .SE(n2627), .CLK(clk), 
        .QN(n2583) );
  SDFFX1_RVT opC10_d4_reg_18_ ( .D(n3424), .SI(1'b0), .SE(n2626), .CLK(clk), 
        .QN(n2581) );
  SDFFX1_RVT opC10_d4_reg_17_ ( .D(n3424), .SI(1'b0), .SE(n2625), .CLK(clk), 
        .QN(n2579) );
  SDFFX1_RVT opC10_d4_reg_16_ ( .D(n3424), .SI(1'b0), .SE(n2624), .CLK(clk), 
        .QN(n2577) );
  SDFFX1_RVT opC10_d4_reg_15_ ( .D(n3424), .SI(1'b0), .SE(n2623), .CLK(clk), 
        .QN(n2575) );
  SDFFX1_RVT opC10_d4_reg_14_ ( .D(n3424), .SI(1'b0), .SE(n2622), .CLK(clk), 
        .QN(n2573) );
  SDFFX1_RVT opC10_d4_reg_13_ ( .D(n3424), .SI(1'b0), .SE(n2621), .CLK(clk), 
        .QN(n2571) );
  SDFFX1_RVT opC10_d4_reg_12_ ( .D(n3424), .SI(1'b0), .SE(n2620), .CLK(clk), 
        .QN(n2569) );
  SDFFX1_RVT opC10_d4_reg_11_ ( .D(n3424), .SI(1'b0), .SE(n2619), .CLK(clk), 
        .QN(n2567) );
  SDFFX1_RVT opC10_d4_reg_10_ ( .D(n3424), .SI(1'b0), .SE(n2618), .CLK(clk), 
        .QN(n2565) );
  SDFFX1_RVT opC10_d4_reg_9_ ( .D(n3424), .SI(1'b0), .SE(n2617), .CLK(clk), 
        .QN(n2563) );
  SDFFX1_RVT opC10_d4_reg_8_ ( .D(n3423), .SI(1'b0), .SE(n2616), .CLK(clk), 
        .QN(n2561) );
  SDFFX1_RVT opC10_d4_reg_7_ ( .D(n3423), .SI(1'b0), .SE(n2615), .CLK(clk), 
        .QN(n2559) );
  SDFFX1_RVT opC10_d4_reg_6_ ( .D(n3423), .SI(1'b0), .SE(n2614), .CLK(clk), 
        .QN(n2557) );
  SDFFX1_RVT opC10_d4_reg_5_ ( .D(n3423), .SI(1'b0), .SE(n2613), .CLK(clk), 
        .QN(n2555) );
  SDFFX1_RVT opC10_d4_reg_4_ ( .D(n3423), .SI(1'b0), .SE(n2612), .CLK(clk), 
        .QN(n2553) );
  SDFFX1_RVT opC10_d4_reg_3_ ( .D(n3423), .SI(1'b0), .SE(n2611), .CLK(clk), 
        .QN(n2551) );
  SDFFX1_RVT opC10_d4_reg_2_ ( .D(n3423), .SI(1'b0), .SE(n2610), .CLK(clk), 
        .QN(n2549) );
  SDFFX1_RVT opC10_d4_reg_1_ ( .D(n3423), .SI(1'b0), .SE(n2609), .CLK(clk), 
        .QN(n2547) );
  SDFFX1_RVT opC10_d4_reg_0_ ( .D(n3423), .SI(1'b0), .SE(n2608), .CLK(clk), 
        .QN(n2545) );
  SDFFX1_RVT opC10_d3_reg_31_ ( .D(n3423), .SI(1'b0), .SE(n2607), .CLK(clk), 
        .QN(n2543) );
  SDFFX1_RVT opC10_d3_reg_30_ ( .D(n3423), .SI(1'b0), .SE(n2605), .CLK(clk), 
        .QN(n2541) );
  SDFFX1_RVT opC10_d3_reg_29_ ( .D(n3423), .SI(1'b0), .SE(n2603), .CLK(clk), 
        .QN(n2539) );
  SDFFX1_RVT opC10_d3_reg_28_ ( .D(n3423), .SI(1'b0), .SE(n2601), .CLK(clk), 
        .QN(n2537) );
  SDFFX1_RVT opC10_d3_reg_27_ ( .D(n3423), .SI(1'b0), .SE(n2599), .CLK(clk), 
        .QN(n2535) );
  SDFFX1_RVT opC10_d3_reg_26_ ( .D(n3422), .SI(1'b0), .SE(n2597), .CLK(clk), 
        .QN(n2533) );
  SDFFX1_RVT opC10_d3_reg_25_ ( .D(n3422), .SI(1'b0), .SE(n2595), .CLK(clk), 
        .QN(n2531) );
  SDFFX1_RVT opC10_d3_reg_24_ ( .D(n3422), .SI(1'b0), .SE(n2593), .CLK(clk), 
        .QN(n2529) );
  SDFFX1_RVT opC10_d3_reg_23_ ( .D(n3422), .SI(1'b0), .SE(n2591), .CLK(clk), 
        .QN(n2527) );
  SDFFX1_RVT opC10_d3_reg_22_ ( .D(n3422), .SI(1'b0), .SE(n2589), .CLK(clk), 
        .QN(n2525) );
  SDFFX1_RVT opC10_d3_reg_21_ ( .D(n3422), .SI(1'b0), .SE(n2587), .CLK(clk), 
        .QN(n2523) );
  SDFFX1_RVT opC10_d3_reg_20_ ( .D(n3422), .SI(1'b0), .SE(n2585), .CLK(clk), 
        .QN(n2521) );
  SDFFX1_RVT opC10_d3_reg_19_ ( .D(n3422), .SI(1'b0), .SE(n2583), .CLK(clk), 
        .QN(n2519) );
  SDFFX1_RVT opC10_d3_reg_18_ ( .D(n3422), .SI(1'b0), .SE(n2581), .CLK(clk), 
        .QN(n2517) );
  SDFFX1_RVT opC10_d3_reg_17_ ( .D(n3422), .SI(1'b0), .SE(n2579), .CLK(clk), 
        .QN(n2515) );
  SDFFX1_RVT opC10_d3_reg_16_ ( .D(n3422), .SI(1'b0), .SE(n2577), .CLK(clk), 
        .QN(n2513) );
  SDFFX1_RVT opC10_d3_reg_15_ ( .D(n3422), .SI(1'b0), .SE(n2575), .CLK(clk), 
        .QN(n2511) );
  SDFFX1_RVT opC10_d3_reg_14_ ( .D(n3421), .SI(1'b0), .SE(n2573), .CLK(clk), 
        .QN(n2509) );
  SDFFX1_RVT opC10_d3_reg_13_ ( .D(n3421), .SI(1'b0), .SE(n2571), .CLK(clk), 
        .QN(n2507) );
  SDFFX1_RVT opC10_d3_reg_12_ ( .D(n3421), .SI(1'b0), .SE(n2569), .CLK(clk), 
        .QN(n2505) );
  SDFFX1_RVT opC10_d3_reg_11_ ( .D(n3421), .SI(1'b0), .SE(n2567), .CLK(clk), 
        .QN(n2503) );
  SDFFX1_RVT opC10_d3_reg_10_ ( .D(n3421), .SI(1'b0), .SE(n2565), .CLK(clk), 
        .QN(n2501) );
  SDFFX1_RVT opC10_d3_reg_9_ ( .D(n3421), .SI(1'b0), .SE(n2563), .CLK(clk), 
        .QN(n2499) );
  SDFFX1_RVT opC10_d3_reg_8_ ( .D(n3421), .SI(1'b0), .SE(n2561), .CLK(clk), 
        .QN(n2497) );
  SDFFX1_RVT opC10_d3_reg_7_ ( .D(n3421), .SI(1'b0), .SE(n2559), .CLK(clk), 
        .QN(n2495) );
  SDFFX1_RVT opC10_d3_reg_6_ ( .D(n3421), .SI(1'b0), .SE(n2557), .CLK(clk), 
        .QN(n2493) );
  SDFFX1_RVT opC10_d3_reg_5_ ( .D(n3421), .SI(1'b0), .SE(n2555), .CLK(clk), 
        .QN(n2491) );
  SDFFX1_RVT opC10_d3_reg_4_ ( .D(n3421), .SI(1'b0), .SE(n2553), .CLK(clk), 
        .QN(n2489) );
  SDFFX1_RVT opC10_d3_reg_3_ ( .D(n3421), .SI(1'b0), .SE(n2551), .CLK(clk), 
        .QN(n2487) );
  SDFFX1_RVT opC10_d3_reg_2_ ( .D(n3421), .SI(1'b0), .SE(n2549), .CLK(clk), 
        .QN(n2485) );
  SDFFX1_RVT opC10_d3_reg_1_ ( .D(n3421), .SI(1'b0), .SE(n2547), .CLK(clk), 
        .QN(n2483) );
  SDFFX1_RVT opC10_d3_reg_0_ ( .D(n3420), .SI(1'b0), .SE(n2545), .CLK(clk), 
        .QN(n2481) );
  SDFFX1_RVT opC10_d2_reg_31_ ( .D(n3420), .SI(1'b0), .SE(n2543), .CLK(clk), 
        .QN(n2479) );
  SDFFX1_RVT opC10_d2_reg_30_ ( .D(n3420), .SI(1'b0), .SE(n2541), .CLK(clk), 
        .QN(n2477) );
  SDFFX1_RVT opC10_d2_reg_29_ ( .D(n3420), .SI(1'b0), .SE(n2539), .CLK(clk), 
        .QN(n2475) );
  SDFFX1_RVT opC10_d2_reg_28_ ( .D(n3420), .SI(1'b0), .SE(n2537), .CLK(clk), 
        .QN(n2473) );
  SDFFX1_RVT opC10_d2_reg_27_ ( .D(n3420), .SI(1'b0), .SE(n2535), .CLK(clk), 
        .QN(n2471) );
  SDFFX1_RVT opC10_d2_reg_26_ ( .D(n3420), .SI(1'b0), .SE(n2533), .CLK(clk), 
        .QN(n2469) );
  SDFFX1_RVT opC10_d2_reg_25_ ( .D(n3420), .SI(1'b0), .SE(n2531), .CLK(clk), 
        .QN(n2467) );
  SDFFX1_RVT opC10_d2_reg_24_ ( .D(n3420), .SI(1'b0), .SE(n2529), .CLK(clk), 
        .QN(n2465) );
  SDFFX1_RVT opC10_d2_reg_23_ ( .D(n3420), .SI(1'b0), .SE(n2527), .CLK(clk), 
        .QN(n2463) );
  SDFFX1_RVT opC10_d2_reg_22_ ( .D(n3420), .SI(1'b0), .SE(n2525), .CLK(clk), 
        .QN(n2461) );
  SDFFX1_RVT opC10_d2_reg_21_ ( .D(n3420), .SI(1'b0), .SE(n2523), .CLK(clk), 
        .QN(n2459) );
  SDFFX1_RVT opC10_d2_reg_20_ ( .D(n3420), .SI(1'b0), .SE(n2521), .CLK(clk), 
        .QN(n2457) );
  SDFFX1_RVT opC10_d2_reg_19_ ( .D(n3420), .SI(1'b0), .SE(n2519), .CLK(clk), 
        .QN(n2455) );
  SDFFX1_RVT opC10_d2_reg_18_ ( .D(n3419), .SI(1'b0), .SE(n2517), .CLK(clk), 
        .QN(n2453) );
  SDFFX1_RVT opC10_d2_reg_17_ ( .D(n3419), .SI(1'b0), .SE(n2515), .CLK(clk), 
        .QN(n2451) );
  SDFFX1_RVT opC10_d2_reg_16_ ( .D(n3419), .SI(1'b0), .SE(n2513), .CLK(clk), 
        .QN(n2449) );
  SDFFX1_RVT opC10_d2_reg_15_ ( .D(n3419), .SI(1'b0), .SE(n2511), .CLK(clk), 
        .QN(n2447) );
  SDFFX1_RVT opC10_d2_reg_14_ ( .D(n3419), .SI(1'b0), .SE(n2509), .CLK(clk), 
        .QN(n2445) );
  SDFFX1_RVT opC10_d2_reg_13_ ( .D(n3419), .SI(1'b0), .SE(n2507), .CLK(clk), 
        .QN(n2443) );
  SDFFX1_RVT opC10_d2_reg_12_ ( .D(n3419), .SI(1'b0), .SE(n2505), .CLK(clk), 
        .QN(n2441) );
  SDFFX1_RVT opC10_d2_reg_11_ ( .D(n3419), .SI(1'b0), .SE(n2503), .CLK(clk), 
        .QN(n2439) );
  SDFFX1_RVT opC10_d2_reg_10_ ( .D(n3419), .SI(1'b0), .SE(n2501), .CLK(clk), 
        .QN(n2437) );
  SDFFX1_RVT opC10_d2_reg_9_ ( .D(n3419), .SI(1'b0), .SE(n2499), .CLK(clk), 
        .QN(n2435) );
  SDFFX1_RVT opC10_d2_reg_8_ ( .D(n3419), .SI(1'b0), .SE(n2497), .CLK(clk), 
        .QN(n2433) );
  SDFFX1_RVT opC10_d2_reg_7_ ( .D(n3419), .SI(1'b0), .SE(n2495), .CLK(clk), 
        .QN(n2431) );
  SDFFX1_RVT opC10_d2_reg_6_ ( .D(n3419), .SI(1'b0), .SE(n2493), .CLK(clk), 
        .QN(n2429) );
  SDFFX1_RVT opC10_d2_reg_5_ ( .D(n3419), .SI(1'b0), .SE(n2491), .CLK(clk), 
        .QN(n2427) );
  SDFFX1_RVT opC10_d2_reg_4_ ( .D(n3418), .SI(1'b0), .SE(n2489), .CLK(clk), 
        .QN(n2425) );
  SDFFX1_RVT opC10_d2_reg_3_ ( .D(n3418), .SI(1'b0), .SE(n2487), .CLK(clk), 
        .QN(n2423) );
  SDFFX1_RVT opC10_d2_reg_2_ ( .D(n3418), .SI(1'b0), .SE(n2485), .CLK(clk), 
        .QN(n2421) );
  SDFFX1_RVT opC10_d2_reg_1_ ( .D(n3418), .SI(1'b0), .SE(n2483), .CLK(clk), 
        .QN(n2419) );
  SDFFX1_RVT opC10_d2_reg_0_ ( .D(n3418), .SI(1'b0), .SE(n2481), .CLK(clk), 
        .QN(n2417) );
  SDFFX1_RVT opC10_d1_reg_31_ ( .D(n3418), .SI(1'b0), .SE(n2479), .CLK(clk), 
        .Q(OpC10[31]) );
  SDFFX1_RVT opC10_d1_reg_30_ ( .D(n3418), .SI(1'b0), .SE(n2477), .CLK(clk), 
        .Q(OpC10[30]) );
  SDFFX1_RVT opC10_d1_reg_29_ ( .D(n3418), .SI(1'b0), .SE(n2475), .CLK(clk), 
        .Q(OpC10[29]) );
  SDFFX1_RVT opC10_d1_reg_28_ ( .D(n3418), .SI(1'b0), .SE(n2473), .CLK(clk), 
        .Q(OpC10[28]) );
  SDFFX1_RVT opC10_d1_reg_27_ ( .D(n3418), .SI(1'b0), .SE(n2471), .CLK(clk), 
        .Q(OpC10[27]) );
  SDFFX1_RVT opC10_d1_reg_26_ ( .D(n3418), .SI(1'b0), .SE(n2469), .CLK(clk), 
        .Q(OpC10[26]) );
  SDFFX1_RVT opC10_d1_reg_25_ ( .D(n3427), .SI(1'b0), .SE(n2467), .CLK(clk), 
        .Q(OpC10[25]) );
  SDFFX1_RVT opC10_d1_reg_24_ ( .D(n3418), .SI(1'b0), .SE(n2465), .CLK(clk), 
        .Q(OpC10[24]) );
  SDFFX1_RVT opC10_d1_reg_23_ ( .D(n3422), .SI(1'b0), .SE(n2463), .CLK(clk), 
        .Q(OpC10[23]) );
  SDFFX1_RVT opC10_d1_reg_22_ ( .D(n3418), .SI(1'b0), .SE(n2461), .CLK(clk), 
        .Q(OpC10[22]) );
  SDFFX1_RVT opC10_d1_reg_21_ ( .D(n3427), .SI(1'b0), .SE(n2459), .CLK(clk), 
        .Q(OpC10[21]) );
  SDFFX1_RVT opC10_d1_reg_20_ ( .D(n3381), .SI(1'b0), .SE(n2457), .CLK(clk), 
        .Q(OpC10[20]) );
  SDFFX1_RVT opC10_d1_reg_19_ ( .D(n3417), .SI(1'b0), .SE(n2455), .CLK(clk), 
        .Q(OpC10[19]) );
  SDFFX1_RVT opC10_d1_reg_18_ ( .D(n3417), .SI(1'b0), .SE(n2453), .CLK(clk), 
        .Q(OpC10[18]) );
  SDFFX1_RVT opC10_d1_reg_17_ ( .D(n3417), .SI(1'b0), .SE(n2451), .CLK(clk), 
        .Q(OpC10[17]) );
  SDFFX1_RVT opC10_d1_reg_16_ ( .D(n3417), .SI(1'b0), .SE(n2449), .CLK(clk), 
        .Q(OpC10[16]) );
  SDFFX1_RVT opC10_d1_reg_15_ ( .D(n3417), .SI(1'b0), .SE(n2447), .CLK(clk), 
        .Q(OpC10[15]) );
  SDFFX1_RVT opC10_d1_reg_14_ ( .D(n3417), .SI(1'b0), .SE(n2445), .CLK(clk), 
        .Q(OpC10[14]) );
  SDFFX1_RVT opC10_d1_reg_13_ ( .D(n3417), .SI(1'b0), .SE(n2443), .CLK(clk), 
        .Q(OpC10[13]) );
  SDFFX1_RVT opC10_d1_reg_12_ ( .D(n3417), .SI(1'b0), .SE(n2441), .CLK(clk), 
        .Q(OpC10[12]) );
  SDFFX1_RVT opC10_d1_reg_11_ ( .D(n3417), .SI(1'b0), .SE(n2439), .CLK(clk), 
        .Q(OpC10[11]) );
  SDFFX1_RVT opC10_d1_reg_10_ ( .D(n3417), .SI(1'b0), .SE(n2437), .CLK(clk), 
        .Q(OpC10[10]) );
  SDFFX1_RVT opC10_d1_reg_9_ ( .D(n3417), .SI(1'b0), .SE(n2435), .CLK(clk), 
        .Q(OpC10[9]) );
  SDFFX1_RVT opC10_d1_reg_8_ ( .D(n3417), .SI(1'b0), .SE(n2433), .CLK(clk), 
        .Q(OpC10[8]) );
  SDFFX1_RVT opC10_d1_reg_7_ ( .D(n3417), .SI(1'b0), .SE(n2431), .CLK(clk), 
        .Q(OpC10[7]) );
  SDFFX1_RVT opC10_d1_reg_6_ ( .D(n3416), .SI(1'b0), .SE(n2429), .CLK(clk), 
        .Q(OpC10[6]) );
  SDFFX1_RVT opC10_d1_reg_5_ ( .D(n3416), .SI(1'b0), .SE(n2427), .CLK(clk), 
        .Q(OpC10[5]) );
  SDFFX1_RVT opC10_d1_reg_4_ ( .D(n3416), .SI(1'b0), .SE(n2425), .CLK(clk), 
        .Q(OpC10[4]) );
  SDFFX1_RVT opC10_d1_reg_3_ ( .D(n3416), .SI(1'b0), .SE(n2423), .CLK(clk), 
        .Q(OpC10[3]) );
  SDFFX1_RVT opC10_d1_reg_2_ ( .D(n3416), .SI(1'b0), .SE(n2421), .CLK(clk), 
        .Q(OpC10[2]) );
  SDFFX1_RVT opC10_d1_reg_1_ ( .D(n3416), .SI(1'b0), .SE(n2419), .CLK(clk), 
        .Q(OpC10[1]) );
  SDFFX1_RVT opC10_d1_reg_0_ ( .D(n3416), .SI(1'b0), .SE(n2417), .CLK(clk), 
        .Q(OpC10[0]) );
  SDFFX1_RVT opC02_d3_reg_31_ ( .D(n3416), .SI(1'b0), .SE(n2383), .CLK(clk), 
        .QN(n2351) );
  SDFFX1_RVT opC02_d3_reg_30_ ( .D(n3416), .SI(1'b0), .SE(n2382), .CLK(clk), 
        .QN(n2349) );
  SDFFX1_RVT opC02_d3_reg_29_ ( .D(n3416), .SI(1'b0), .SE(n2381), .CLK(clk), 
        .QN(n2347) );
  SDFFX1_RVT opC02_d3_reg_28_ ( .D(n3416), .SI(1'b0), .SE(n2380), .CLK(clk), 
        .QN(n2345) );
  SDFFX1_RVT opC02_d3_reg_27_ ( .D(n3416), .SI(1'b0), .SE(n2379), .CLK(clk), 
        .QN(n2343) );
  SDFFX1_RVT opC02_d3_reg_26_ ( .D(n3416), .SI(1'b0), .SE(n2378), .CLK(clk), 
        .QN(n2341) );
  SDFFX1_RVT opC02_d3_reg_25_ ( .D(n3416), .SI(1'b0), .SE(n2377), .CLK(clk), 
        .QN(n2339) );
  SDFFX1_RVT opC02_d3_reg_24_ ( .D(n3415), .SI(1'b0), .SE(n2376), .CLK(clk), 
        .QN(n2337) );
  SDFFX1_RVT opC02_d3_reg_23_ ( .D(n3415), .SI(1'b0), .SE(n2375), .CLK(clk), 
        .QN(n2335) );
  SDFFX1_RVT opC02_d3_reg_22_ ( .D(n3415), .SI(1'b0), .SE(n2374), .CLK(clk), 
        .QN(n2333) );
  SDFFX1_RVT opC02_d3_reg_21_ ( .D(n3415), .SI(1'b0), .SE(n2373), .CLK(clk), 
        .QN(n2331) );
  SDFFX1_RVT opC02_d3_reg_20_ ( .D(n3415), .SI(1'b0), .SE(n2372), .CLK(clk), 
        .QN(n2329) );
  SDFFX1_RVT opC02_d3_reg_19_ ( .D(n3415), .SI(1'b0), .SE(n2371), .CLK(clk), 
        .QN(n2327) );
  SDFFX1_RVT opC02_d3_reg_18_ ( .D(n3415), .SI(1'b0), .SE(n2370), .CLK(clk), 
        .QN(n2325) );
  SDFFX1_RVT opC02_d3_reg_17_ ( .D(n3415), .SI(1'b0), .SE(n2369), .CLK(clk), 
        .QN(n2323) );
  SDFFX1_RVT opC02_d3_reg_16_ ( .D(n3415), .SI(1'b0), .SE(n2368), .CLK(clk), 
        .QN(n2321) );
  SDFFX1_RVT opC02_d3_reg_15_ ( .D(n3415), .SI(1'b0), .SE(n2367), .CLK(clk), 
        .QN(n2319) );
  SDFFX1_RVT opC02_d3_reg_14_ ( .D(n3415), .SI(1'b0), .SE(n2366), .CLK(clk), 
        .QN(n2317) );
  SDFFX1_RVT opC02_d3_reg_13_ ( .D(n3415), .SI(1'b0), .SE(n2365), .CLK(clk), 
        .QN(n2315) );
  SDFFX1_RVT opC02_d3_reg_12_ ( .D(n3415), .SI(1'b0), .SE(n2364), .CLK(clk), 
        .QN(n2313) );
  SDFFX1_RVT opC02_d3_reg_11_ ( .D(n3415), .SI(1'b0), .SE(n2363), .CLK(clk), 
        .QN(n2311) );
  SDFFX1_RVT opC02_d3_reg_10_ ( .D(n3414), .SI(1'b0), .SE(n2362), .CLK(clk), 
        .QN(n2309) );
  SDFFX1_RVT opC02_d3_reg_9_ ( .D(n3414), .SI(1'b0), .SE(n2361), .CLK(clk), 
        .QN(n2307) );
  SDFFX1_RVT opC02_d3_reg_8_ ( .D(n3414), .SI(1'b0), .SE(n2360), .CLK(clk), 
        .QN(n2305) );
  SDFFX1_RVT opC02_d3_reg_7_ ( .D(n3414), .SI(1'b0), .SE(n2359), .CLK(clk), 
        .QN(n2303) );
  SDFFX1_RVT opC02_d3_reg_6_ ( .D(n3414), .SI(1'b0), .SE(n2358), .CLK(clk), 
        .QN(n2301) );
  SDFFX1_RVT opC02_d3_reg_5_ ( .D(n3414), .SI(1'b0), .SE(n2357), .CLK(clk), 
        .QN(n2299) );
  SDFFX1_RVT opC02_d3_reg_4_ ( .D(n3414), .SI(1'b0), .SE(n2356), .CLK(clk), 
        .QN(n2297) );
  SDFFX1_RVT opC02_d3_reg_3_ ( .D(n3414), .SI(1'b0), .SE(n2355), .CLK(clk), 
        .QN(n2295) );
  SDFFX1_RVT opC02_d3_reg_2_ ( .D(n3414), .SI(1'b0), .SE(n2354), .CLK(clk), 
        .QN(n2293) );
  SDFFX1_RVT opC02_d3_reg_1_ ( .D(n3414), .SI(1'b0), .SE(n2353), .CLK(clk), 
        .QN(n2291) );
  SDFFX1_RVT opC02_d3_reg_0_ ( .D(n3414), .SI(1'b0), .SE(n2352), .CLK(clk), 
        .QN(n2289) );
  SDFFX1_RVT opC02_d2_reg_31_ ( .D(n3414), .SI(1'b0), .SE(n2351), .CLK(clk), 
        .QN(n2287) );
  SDFFX1_RVT opC02_d2_reg_30_ ( .D(n3414), .SI(1'b0), .SE(n2349), .CLK(clk), 
        .QN(n2285) );
  SDFFX1_RVT opC02_d2_reg_29_ ( .D(n3414), .SI(1'b0), .SE(n2347), .CLK(clk), 
        .QN(n2283) );
  SDFFX1_RVT opC02_d2_reg_28_ ( .D(n3413), .SI(1'b0), .SE(n2345), .CLK(clk), 
        .QN(n2281) );
  SDFFX1_RVT opC02_d2_reg_27_ ( .D(n3413), .SI(1'b0), .SE(n2343), .CLK(clk), 
        .QN(n2279) );
  SDFFX1_RVT opC02_d2_reg_26_ ( .D(n3413), .SI(1'b0), .SE(n2341), .CLK(clk), 
        .QN(n2277) );
  SDFFX1_RVT opC02_d2_reg_25_ ( .D(n3413), .SI(1'b0), .SE(n2339), .CLK(clk), 
        .QN(n2275) );
  SDFFX1_RVT opC02_d2_reg_24_ ( .D(n3413), .SI(1'b0), .SE(n2337), .CLK(clk), 
        .QN(n2273) );
  SDFFX1_RVT opC02_d2_reg_23_ ( .D(n3413), .SI(1'b0), .SE(n2335), .CLK(clk), 
        .QN(n2271) );
  SDFFX1_RVT opC02_d2_reg_22_ ( .D(n3413), .SI(1'b0), .SE(n2333), .CLK(clk), 
        .QN(n2269) );
  SDFFX1_RVT opC02_d2_reg_21_ ( .D(n3413), .SI(1'b0), .SE(n2331), .CLK(clk), 
        .QN(n2267) );
  SDFFX1_RVT opC02_d2_reg_20_ ( .D(n3413), .SI(1'b0), .SE(n2329), .CLK(clk), 
        .QN(n2265) );
  SDFFX1_RVT opC02_d2_reg_19_ ( .D(n3413), .SI(1'b0), .SE(n2327), .CLK(clk), 
        .QN(n2263) );
  SDFFX1_RVT opC02_d2_reg_18_ ( .D(n3413), .SI(1'b0), .SE(n2325), .CLK(clk), 
        .QN(n2261) );
  SDFFX1_RVT opC02_d2_reg_17_ ( .D(n3413), .SI(1'b0), .SE(n2323), .CLK(clk), 
        .QN(n2259) );
  SDFFX1_RVT opC02_d2_reg_16_ ( .D(n3412), .SI(1'b0), .SE(n2321), .CLK(clk), 
        .QN(n2257) );
  SDFFX1_RVT opC02_d2_reg_15_ ( .D(n3412), .SI(1'b0), .SE(n2319), .CLK(clk), 
        .QN(n2255) );
  SDFFX1_RVT opC02_d2_reg_14_ ( .D(n3412), .SI(1'b0), .SE(n2317), .CLK(clk), 
        .QN(n2253) );
  SDFFX1_RVT opC02_d2_reg_13_ ( .D(n3412), .SI(1'b0), .SE(n2315), .CLK(clk), 
        .QN(n2251) );
  SDFFX1_RVT opC02_d2_reg_12_ ( .D(n3412), .SI(1'b0), .SE(n2313), .CLK(clk), 
        .QN(n2249) );
  SDFFX1_RVT opC02_d2_reg_11_ ( .D(n3412), .SI(1'b0), .SE(n2311), .CLK(clk), 
        .QN(n2247) );
  SDFFX1_RVT opC02_d2_reg_10_ ( .D(n3412), .SI(1'b0), .SE(n2309), .CLK(clk), 
        .QN(n2245) );
  SDFFX1_RVT opC02_d2_reg_9_ ( .D(n3412), .SI(1'b0), .SE(n2307), .CLK(clk), 
        .QN(n2243) );
  SDFFX1_RVT opC02_d2_reg_8_ ( .D(n3412), .SI(1'b0), .SE(n2305), .CLK(clk), 
        .QN(n2241) );
  SDFFX1_RVT opC02_d2_reg_7_ ( .D(n3412), .SI(1'b0), .SE(n2303), .CLK(clk), 
        .QN(n2239) );
  SDFFX1_RVT opC02_d2_reg_6_ ( .D(n3412), .SI(1'b0), .SE(n2301), .CLK(clk), 
        .QN(n2237) );
  SDFFX1_RVT opC02_d2_reg_5_ ( .D(n3412), .SI(1'b0), .SE(n2299), .CLK(clk), 
        .QN(n2235) );
  SDFFX1_RVT opC02_d2_reg_4_ ( .D(n3412), .SI(1'b0), .SE(n2297), .CLK(clk), 
        .QN(n2233) );
  SDFFX1_RVT opC02_d2_reg_3_ ( .D(n3412), .SI(1'b0), .SE(n2295), .CLK(clk), 
        .QN(n2231) );
  SDFFX1_RVT opC02_d2_reg_2_ ( .D(n3411), .SI(1'b0), .SE(n2293), .CLK(clk), 
        .QN(n2229) );
  SDFFX1_RVT opC02_d2_reg_1_ ( .D(n3411), .SI(1'b0), .SE(n2291), .CLK(clk), 
        .QN(n2227) );
  SDFFX1_RVT opC02_d2_reg_0_ ( .D(n3411), .SI(1'b0), .SE(n2289), .CLK(clk), 
        .QN(n2225) );
  SDFFX1_RVT opC02_d1_reg_31_ ( .D(n3411), .SI(1'b0), .SE(n2287), .CLK(clk), 
        .Q(OpC02[31]) );
  SDFFX1_RVT opC02_d1_reg_30_ ( .D(n3411), .SI(1'b0), .SE(n2285), .CLK(clk), 
        .Q(OpC02[30]) );
  SDFFX1_RVT opC02_d1_reg_29_ ( .D(n3411), .SI(1'b0), .SE(n2283), .CLK(clk), 
        .Q(OpC02[29]) );
  SDFFX1_RVT opC02_d1_reg_28_ ( .D(n3411), .SI(1'b0), .SE(n2281), .CLK(clk), 
        .Q(OpC02[28]) );
  SDFFX1_RVT opC02_d1_reg_27_ ( .D(n3411), .SI(1'b0), .SE(n2279), .CLK(clk), 
        .Q(OpC02[27]) );
  SDFFX1_RVT opC02_d1_reg_26_ ( .D(n3411), .SI(1'b0), .SE(n2277), .CLK(clk), 
        .Q(OpC02[26]) );
  SDFFX1_RVT opC02_d1_reg_25_ ( .D(n3411), .SI(1'b0), .SE(n2275), .CLK(clk), 
        .Q(OpC02[25]) );
  SDFFX1_RVT opC02_d1_reg_24_ ( .D(n3411), .SI(1'b0), .SE(n2273), .CLK(clk), 
        .Q(OpC02[24]) );
  SDFFX1_RVT opC02_d1_reg_23_ ( .D(n3411), .SI(1'b0), .SE(n2271), .CLK(clk), 
        .Q(OpC02[23]) );
  SDFFX1_RVT opC02_d1_reg_22_ ( .D(n3411), .SI(1'b0), .SE(n2269), .CLK(clk), 
        .Q(OpC02[22]) );
  SDFFX1_RVT opC02_d1_reg_21_ ( .D(n3411), .SI(1'b0), .SE(n2267), .CLK(clk), 
        .Q(OpC02[21]) );
  SDFFX1_RVT opC02_d1_reg_20_ ( .D(n3410), .SI(1'b0), .SE(n2265), .CLK(clk), 
        .Q(OpC02[20]) );
  SDFFX1_RVT opC02_d1_reg_19_ ( .D(n3410), .SI(1'b0), .SE(n2263), .CLK(clk), 
        .Q(OpC02[19]) );
  SDFFX1_RVT opC02_d1_reg_18_ ( .D(n3410), .SI(1'b0), .SE(n2261), .CLK(clk), 
        .Q(OpC02[18]) );
  SDFFX1_RVT opC02_d1_reg_17_ ( .D(n3410), .SI(1'b0), .SE(n2259), .CLK(clk), 
        .Q(OpC02[17]) );
  SDFFX1_RVT opC02_d1_reg_16_ ( .D(n3410), .SI(1'b0), .SE(n2257), .CLK(clk), 
        .Q(OpC02[16]) );
  SDFFX1_RVT opC02_d1_reg_15_ ( .D(n3410), .SI(1'b0), .SE(n2255), .CLK(clk), 
        .Q(OpC02[15]) );
  SDFFX1_RVT opC02_d1_reg_14_ ( .D(n3410), .SI(1'b0), .SE(n2253), .CLK(clk), 
        .Q(OpC02[14]) );
  SDFFX1_RVT opC02_d1_reg_13_ ( .D(n3410), .SI(1'b0), .SE(n2251), .CLK(clk), 
        .Q(OpC02[13]) );
  SDFFX1_RVT opC02_d1_reg_12_ ( .D(n3410), .SI(1'b0), .SE(n2249), .CLK(clk), 
        .Q(OpC02[12]) );
  SDFFX1_RVT opC02_d1_reg_11_ ( .D(n3410), .SI(1'b0), .SE(n2247), .CLK(clk), 
        .Q(OpC02[11]) );
  SDFFX1_RVT opC02_d1_reg_10_ ( .D(n3410), .SI(1'b0), .SE(n2245), .CLK(clk), 
        .Q(OpC02[10]) );
  SDFFX1_RVT opC02_d1_reg_9_ ( .D(n3410), .SI(1'b0), .SE(n2243), .CLK(clk), 
        .Q(OpC02[9]) );
  SDFFX1_RVT opC02_d1_reg_8_ ( .D(n3410), .SI(1'b0), .SE(n2241), .CLK(clk), 
        .Q(OpC02[8]) );
  SDFFX1_RVT opC02_d1_reg_7_ ( .D(n3410), .SI(1'b0), .SE(n2239), .CLK(clk), 
        .Q(OpC02[7]) );
  SDFFX1_RVT opC02_d1_reg_6_ ( .D(n3409), .SI(1'b0), .SE(n2237), .CLK(clk), 
        .Q(OpC02[6]) );
  SDFFX1_RVT opC02_d1_reg_5_ ( .D(n3409), .SI(1'b0), .SE(n2235), .CLK(clk), 
        .Q(OpC02[5]) );
  SDFFX1_RVT opC02_d1_reg_4_ ( .D(n3409), .SI(1'b0), .SE(n2233), .CLK(clk), 
        .Q(OpC02[4]) );
  SDFFX1_RVT opC02_d1_reg_3_ ( .D(n3409), .SI(1'b0), .SE(n2231), .CLK(clk), 
        .Q(OpC02[3]) );
  SDFFX1_RVT opC02_d1_reg_2_ ( .D(n3409), .SI(1'b0), .SE(n2229), .CLK(clk), 
        .Q(OpC02[2]) );
  SDFFX1_RVT opC02_d1_reg_1_ ( .D(n3409), .SI(1'b0), .SE(n2227), .CLK(clk), 
        .Q(OpC02[1]) );
  SDFFX1_RVT opC02_d1_reg_0_ ( .D(n3409), .SI(1'b0), .SE(n2225), .CLK(clk), 
        .Q(OpC02[0]) );
  SDFFX1_RVT opC11_d3_reg_31_ ( .D(n3409), .SI(1'b0), .SE(n2191), .CLK(clk), 
        .QN(n2159) );
  SDFFX1_RVT opC11_d3_reg_30_ ( .D(n3409), .SI(1'b0), .SE(n2190), .CLK(clk), 
        .QN(n2157) );
  SDFFX1_RVT opC11_d3_reg_29_ ( .D(n3409), .SI(1'b0), .SE(n2189), .CLK(clk), 
        .QN(n2155) );
  SDFFX1_RVT opC11_d3_reg_28_ ( .D(n3409), .SI(1'b0), .SE(n2188), .CLK(clk), 
        .QN(n2153) );
  SDFFX1_RVT opC11_d3_reg_27_ ( .D(n3409), .SI(1'b0), .SE(n2187), .CLK(clk), 
        .QN(n2151) );
  SDFFX1_RVT opC11_d3_reg_26_ ( .D(n3409), .SI(1'b0), .SE(n2186), .CLK(clk), 
        .QN(n2149) );
  SDFFX1_RVT opC11_d3_reg_25_ ( .D(n3409), .SI(1'b0), .SE(n2185), .CLK(clk), 
        .QN(n2147) );
  SDFFX1_RVT opC11_d3_reg_24_ ( .D(n3408), .SI(1'b0), .SE(n2184), .CLK(clk), 
        .QN(n2145) );
  SDFFX1_RVT opC11_d3_reg_23_ ( .D(n3408), .SI(1'b0), .SE(n2183), .CLK(clk), 
        .QN(n2143) );
  SDFFX1_RVT opC11_d3_reg_22_ ( .D(n3408), .SI(1'b0), .SE(n2182), .CLK(clk), 
        .QN(n2141) );
  SDFFX1_RVT opC11_d3_reg_21_ ( .D(n3408), .SI(1'b0), .SE(n2181), .CLK(clk), 
        .QN(n2139) );
  SDFFX1_RVT opC11_d3_reg_20_ ( .D(n3408), .SI(1'b0), .SE(n2180), .CLK(clk), 
        .QN(n2137) );
  SDFFX1_RVT opC11_d3_reg_19_ ( .D(n3413), .SI(1'b0), .SE(n2179), .CLK(clk), 
        .QN(n2135) );
  SDFFX1_RVT opC11_d3_reg_18_ ( .D(n3427), .SI(1'b0), .SE(n2178), .CLK(clk), 
        .QN(n2133) );
  SDFFX1_RVT opC11_d3_reg_17_ ( .D(n3417), .SI(1'b0), .SE(n2177), .CLK(clk), 
        .QN(n2131) );
  SDFFX1_RVT opC11_d3_reg_16_ ( .D(n3394), .SI(1'b0), .SE(n2176), .CLK(clk), 
        .QN(n2129) );
  SDFFX1_RVT opC11_d3_reg_15_ ( .D(n3408), .SI(1'b0), .SE(n2175), .CLK(clk), 
        .QN(n2127) );
  SDFFX1_RVT opC11_d3_reg_14_ ( .D(n3408), .SI(1'b0), .SE(n2174), .CLK(clk), 
        .QN(n2125) );
  SDFFX1_RVT opC11_d3_reg_13_ ( .D(n3408), .SI(1'b0), .SE(n2173), .CLK(clk), 
        .QN(n2123) );
  SDFFX1_RVT opC11_d3_reg_12_ ( .D(n3408), .SI(1'b0), .SE(n2172), .CLK(clk), 
        .QN(n2121) );
  SDFFX1_RVT opC11_d3_reg_11_ ( .D(n3408), .SI(1'b0), .SE(n2171), .CLK(clk), 
        .QN(n2119) );
  SDFFX1_RVT opC11_d3_reg_10_ ( .D(n3408), .SI(1'b0), .SE(n2170), .CLK(clk), 
        .QN(n2117) );
  SDFFX1_RVT opC11_d3_reg_9_ ( .D(n3408), .SI(1'b0), .SE(n2169), .CLK(clk), 
        .QN(n2115) );
  SDFFX1_RVT opC11_d3_reg_8_ ( .D(n3408), .SI(1'b0), .SE(n2168), .CLK(clk), 
        .QN(n2113) );
  SDFFX1_RVT opC11_d3_reg_7_ ( .D(n3407), .SI(1'b0), .SE(n2167), .CLK(clk), 
        .QN(n2111) );
  SDFFX1_RVT opC11_d3_reg_6_ ( .D(n3407), .SI(1'b0), .SE(n2166), .CLK(clk), 
        .Q(opC11_d3_6_) );
  SDFFX1_RVT opC11_d3_reg_5_ ( .D(n3407), .SI(1'b0), .SE(n2165), .CLK(clk), 
        .QN(n2108) );
  SDFFX1_RVT opC11_d3_reg_4_ ( .D(n3407), .SI(1'b0), .SE(n2164), .CLK(clk), 
        .QN(n2106) );
  SDFFX1_RVT opC11_d3_reg_3_ ( .D(n3407), .SI(1'b0), .SE(n2163), .CLK(clk), 
        .QN(n2104) );
  SDFFX1_RVT opC11_d3_reg_2_ ( .D(n3407), .SI(1'b0), .SE(n2162), .CLK(clk), 
        .QN(n2102) );
  SDFFX1_RVT opC11_d3_reg_1_ ( .D(n3407), .SI(1'b0), .SE(n2161), .CLK(clk), 
        .QN(n2100) );
  SDFFX1_RVT opC11_d3_reg_0_ ( .D(n3407), .SI(1'b0), .SE(n2160), .CLK(clk), 
        .QN(n2098) );
  SDFFX1_RVT opC11_d2_reg_31_ ( .D(n3407), .SI(1'b0), .SE(n2159), .CLK(clk), 
        .QN(n2096) );
  SDFFX1_RVT opC11_d2_reg_30_ ( .D(n3407), .SI(1'b0), .SE(n2157), .CLK(clk), 
        .QN(n2094) );
  SDFFX1_RVT opC11_d2_reg_29_ ( .D(n3407), .SI(1'b0), .SE(n2155), .CLK(clk), 
        .QN(n2092) );
  SDFFX1_RVT opC11_d2_reg_28_ ( .D(n3407), .SI(1'b0), .SE(n2153), .CLK(clk), 
        .QN(n2090) );
  SDFFX1_RVT opC11_d2_reg_27_ ( .D(n3407), .SI(1'b0), .SE(n2151), .CLK(clk), 
        .QN(n2088) );
  SDFFX1_RVT opC11_d2_reg_26_ ( .D(n3407), .SI(1'b0), .SE(n2149), .CLK(clk), 
        .QN(n2086) );
  SDFFX1_RVT opC11_d2_reg_25_ ( .D(n3406), .SI(1'b0), .SE(n2147), .CLK(clk), 
        .QN(n2084) );
  SDFFX1_RVT opC11_d2_reg_24_ ( .D(n3406), .SI(1'b0), .SE(n2145), .CLK(clk), 
        .QN(n2082) );
  SDFFX1_RVT opC11_d2_reg_23_ ( .D(n3406), .SI(1'b0), .SE(n2143), .CLK(clk), 
        .QN(n2080) );
  SDFFX1_RVT opC11_d2_reg_22_ ( .D(n3406), .SI(1'b0), .SE(n2141), .CLK(clk), 
        .QN(n2078) );
  SDFFX1_RVT opC11_d2_reg_21_ ( .D(n3406), .SI(1'b0), .SE(n2139), .CLK(clk), 
        .QN(n2076) );
  SDFFX1_RVT opC11_d2_reg_20_ ( .D(n3406), .SI(1'b0), .SE(n2137), .CLK(clk), 
        .QN(n2074) );
  SDFFX1_RVT opC11_d2_reg_19_ ( .D(n3406), .SI(1'b0), .SE(n2135), .CLK(clk), 
        .QN(n2072) );
  SDFFX1_RVT opC11_d2_reg_18_ ( .D(n3406), .SI(1'b0), .SE(n2133), .CLK(clk), 
        .QN(n2070) );
  SDFFX1_RVT opC11_d2_reg_17_ ( .D(n3406), .SI(1'b0), .SE(n2131), .CLK(clk), 
        .QN(n2068) );
  SDFFX1_RVT opC11_d2_reg_16_ ( .D(n3406), .SI(1'b0), .SE(n2129), .CLK(clk), 
        .QN(n2066) );
  SDFFX1_RVT opC11_d2_reg_15_ ( .D(n3406), .SI(1'b0), .SE(n2127), .CLK(clk), 
        .QN(n2064) );
  SDFFX1_RVT opC11_d2_reg_14_ ( .D(n3406), .SI(1'b0), .SE(n2125), .CLK(clk), 
        .QN(n2062) );
  SDFFX1_RVT opC11_d2_reg_13_ ( .D(n3406), .SI(1'b0), .SE(n2123), .CLK(clk), 
        .QN(n2060) );
  SDFFX1_RVT opC11_d2_reg_12_ ( .D(n3406), .SI(1'b0), .SE(n2121), .CLK(clk), 
        .QN(n2058) );
  SDFFX1_RVT opC11_d2_reg_11_ ( .D(n3405), .SI(1'b0), .SE(n2119), .CLK(clk), 
        .QN(n2056) );
  SDFFX1_RVT opC11_d2_reg_10_ ( .D(n3405), .SI(1'b0), .SE(n2117), .CLK(clk), 
        .QN(n2054) );
  SDFFX1_RVT opC11_d2_reg_9_ ( .D(n3405), .SI(1'b0), .SE(n2115), .CLK(clk), 
        .QN(n2052) );
  SDFFX1_RVT opC11_d2_reg_8_ ( .D(n3405), .SI(1'b0), .SE(n2113), .CLK(clk), 
        .QN(n2050) );
  SDFFX1_RVT opC11_d2_reg_7_ ( .D(n3405), .SI(1'b0), .SE(n2111), .CLK(clk), 
        .QN(n2048) );
  SDFFX1_RVT opC11_d2_reg_5_ ( .D(n3405), .SI(1'b0), .SE(n2108), .CLK(clk), 
        .QN(n2045) );
  SDFFX1_RVT opC11_d2_reg_4_ ( .D(n3405), .SI(1'b0), .SE(n2106), .CLK(clk), 
        .QN(n2043) );
  SDFFX1_RVT opC11_d2_reg_3_ ( .D(n3405), .SI(1'b0), .SE(n2104), .CLK(clk), 
        .QN(n2041) );
  SDFFX1_RVT opC11_d2_reg_2_ ( .D(n3405), .SI(1'b0), .SE(n2102), .CLK(clk), 
        .QN(n2039) );
  SDFFX1_RVT opC11_d2_reg_1_ ( .D(n3405), .SI(1'b0), .SE(n2100), .CLK(clk), 
        .QN(n2037) );
  SDFFX1_RVT opC11_d2_reg_0_ ( .D(n3405), .SI(1'b0), .SE(n2098), .CLK(clk), 
        .QN(n2035) );
  SDFFX1_RVT opC11_d1_reg_31_ ( .D(n3405), .SI(1'b0), .SE(n2096), .CLK(clk), 
        .Q(OpC11[31]) );
  SDFFX1_RVT opC11_d1_reg_30_ ( .D(n3405), .SI(1'b0), .SE(n2094), .CLK(clk), 
        .Q(OpC11[30]) );
  SDFFX1_RVT opC11_d1_reg_29_ ( .D(n3405), .SI(1'b0), .SE(n2092), .CLK(clk), 
        .Q(OpC11[29]) );
  SDFFX1_RVT opC11_d1_reg_28_ ( .D(n3404), .SI(1'b0), .SE(n2090), .CLK(clk), 
        .Q(OpC11[28]) );
  SDFFX1_RVT opC11_d1_reg_27_ ( .D(n3404), .SI(1'b0), .SE(n2088), .CLK(clk), 
        .Q(OpC11[27]) );
  SDFFX1_RVT opC11_d1_reg_26_ ( .D(n3404), .SI(1'b0), .SE(n2086), .CLK(clk), 
        .Q(OpC11[26]) );
  SDFFX1_RVT opC11_d1_reg_25_ ( .D(n3404), .SI(1'b0), .SE(n2084), .CLK(clk), 
        .Q(OpC11[25]) );
  SDFFX1_RVT opC11_d1_reg_24_ ( .D(n3404), .SI(1'b0), .SE(n2082), .CLK(clk), 
        .Q(OpC11[24]) );
  SDFFX1_RVT opC11_d1_reg_23_ ( .D(n3404), .SI(1'b0), .SE(n2080), .CLK(clk), 
        .Q(OpC11[23]) );
  SDFFX1_RVT opC11_d1_reg_22_ ( .D(n3404), .SI(1'b0), .SE(n2078), .CLK(clk), 
        .Q(OpC11[22]) );
  SDFFX1_RVT opC11_d1_reg_21_ ( .D(n3404), .SI(1'b0), .SE(n2076), .CLK(clk), 
        .Q(OpC11[21]) );
  SDFFX1_RVT opC11_d1_reg_20_ ( .D(n3404), .SI(1'b0), .SE(n2074), .CLK(clk), 
        .Q(OpC11[20]) );
  SDFFX1_RVT opC11_d1_reg_19_ ( .D(n3404), .SI(1'b0), .SE(n2072), .CLK(clk), 
        .Q(OpC11[19]) );
  SDFFX1_RVT opC11_d1_reg_18_ ( .D(n3404), .SI(1'b0), .SE(n2070), .CLK(clk), 
        .Q(OpC11[18]) );
  SDFFX1_RVT opC11_d1_reg_17_ ( .D(n3404), .SI(1'b0), .SE(n2068), .CLK(clk), 
        .Q(OpC11[17]) );
  SDFFX1_RVT opC11_d1_reg_16_ ( .D(n3404), .SI(1'b0), .SE(n2066), .CLK(clk), 
        .Q(OpC11[16]) );
  SDFFX1_RVT opC11_d1_reg_15_ ( .D(n3404), .SI(1'b0), .SE(n2064), .CLK(clk), 
        .Q(OpC11[15]) );
  SDFFX1_RVT opC11_d1_reg_14_ ( .D(n3403), .SI(1'b0), .SE(n2062), .CLK(clk), 
        .Q(OpC11[14]) );
  SDFFX1_RVT opC11_d1_reg_13_ ( .D(n3403), .SI(1'b0), .SE(n2060), .CLK(clk), 
        .Q(OpC11[13]) );
  SDFFX1_RVT opC11_d1_reg_12_ ( .D(n3403), .SI(1'b0), .SE(n2058), .CLK(clk), 
        .Q(OpC11[12]) );
  SDFFX1_RVT opC11_d1_reg_11_ ( .D(n3403), .SI(1'b0), .SE(n2056), .CLK(clk), 
        .Q(OpC11[11]) );
  SDFFX1_RVT opC11_d1_reg_10_ ( .D(n3403), .SI(1'b0), .SE(n2054), .CLK(clk), 
        .Q(OpC11[10]) );
  SDFFX1_RVT opC11_d1_reg_9_ ( .D(n3403), .SI(1'b0), .SE(n2052), .CLK(clk), 
        .Q(OpC11[9]) );
  SDFFX1_RVT opC11_d1_reg_8_ ( .D(n3403), .SI(1'b0), .SE(n2050), .CLK(clk), 
        .Q(OpC11[8]) );
  SDFFX1_RVT opC11_d1_reg_7_ ( .D(n3403), .SI(1'b0), .SE(n2048), .CLK(clk), 
        .Q(OpC11[7]) );
  SDFFX1_RVT opC11_d1_reg_6_ ( .D(n3403), .SI(1'b0), .SE(n2046), .CLK(clk), 
        .Q(OpC11[6]) );
  SDFFX1_RVT opC11_d1_reg_5_ ( .D(n3403), .SI(1'b0), .SE(n2045), .CLK(clk), 
        .Q(OpC11[5]) );
  SDFFX1_RVT opC11_d1_reg_4_ ( .D(n3403), .SI(1'b0), .SE(n2043), .CLK(clk), 
        .Q(OpC11[4]) );
  SDFFX1_RVT opC11_d1_reg_3_ ( .D(n3403), .SI(1'b0), .SE(n2041), .CLK(clk), 
        .Q(OpC11[3]) );
  SDFFX1_RVT opC11_d1_reg_2_ ( .D(n3402), .SI(1'b0), .SE(n2039), .CLK(clk), 
        .Q(OpC11[2]) );
  SDFFX1_RVT opC11_d1_reg_1_ ( .D(n3402), .SI(1'b0), .SE(n2037), .CLK(clk), 
        .Q(OpC11[1]) );
  SDFFX1_RVT opC11_d1_reg_0_ ( .D(n3402), .SI(1'b0), .SE(n2035), .CLK(clk), 
        .Q(OpC11[0]) );
  SDFFX1_RVT opC20_d3_reg_31_ ( .D(n3402), .SI(1'b0), .SE(n2001), .CLK(clk), 
        .QN(n1969) );
  SDFFX1_RVT opC20_d3_reg_30_ ( .D(n3402), .SI(1'b0), .SE(n2000), .CLK(clk), 
        .QN(n1967) );
  SDFFX1_RVT opC20_d3_reg_29_ ( .D(n3402), .SI(1'b0), .SE(n1999), .CLK(clk), 
        .QN(n1965) );
  SDFFX1_RVT opC20_d3_reg_28_ ( .D(n3402), .SI(1'b0), .SE(n1998), .CLK(clk), 
        .QN(n1963) );
  SDFFX1_RVT opC20_d3_reg_27_ ( .D(n3402), .SI(1'b0), .SE(n1997), .CLK(clk), 
        .QN(n1961) );
  SDFFX1_RVT opC20_d3_reg_26_ ( .D(n3402), .SI(1'b0), .SE(n1996), .CLK(clk), 
        .QN(n1959) );
  SDFFX1_RVT opC20_d3_reg_25_ ( .D(n3402), .SI(1'b0), .SE(n1995), .CLK(clk), 
        .QN(n1957) );
  SDFFX1_RVT opC20_d3_reg_24_ ( .D(n3402), .SI(1'b0), .SE(n1994), .CLK(clk), 
        .QN(n1955) );
  SDFFX1_RVT opC20_d3_reg_23_ ( .D(n3402), .SI(1'b0), .SE(n1993), .CLK(clk), 
        .QN(n1953) );
  SDFFX1_RVT opC20_d3_reg_22_ ( .D(n3402), .SI(1'b0), .SE(n1992), .CLK(clk), 
        .QN(n1951) );
  SDFFX1_RVT opC20_d3_reg_21_ ( .D(n3402), .SI(1'b0), .SE(n1991), .CLK(clk), 
        .QN(n1949) );
  SDFFX1_RVT opC20_d3_reg_20_ ( .D(n3401), .SI(1'b0), .SE(n1990), .CLK(clk), 
        .QN(n1947) );
  SDFFX1_RVT opC20_d3_reg_19_ ( .D(n3401), .SI(1'b0), .SE(n1989), .CLK(clk), 
        .QN(n1945) );
  SDFFX1_RVT opC20_d3_reg_18_ ( .D(n3401), .SI(1'b0), .SE(n1988), .CLK(clk), 
        .QN(n1943) );
  SDFFX1_RVT opC20_d3_reg_17_ ( .D(n3401), .SI(1'b0), .SE(n1987), .CLK(clk), 
        .QN(n1941) );
  SDFFX1_RVT opC20_d3_reg_16_ ( .D(n3401), .SI(1'b0), .SE(n1986), .CLK(clk), 
        .QN(n1939) );
  SDFFX1_RVT opC20_d3_reg_15_ ( .D(n3401), .SI(1'b0), .SE(n1985), .CLK(clk), 
        .QN(n1937) );
  SDFFX1_RVT opC20_d3_reg_14_ ( .D(n3401), .SI(1'b0), .SE(n1984), .CLK(clk), 
        .QN(n1935) );
  SDFFX1_RVT opC20_d3_reg_13_ ( .D(n3401), .SI(1'b0), .SE(n1983), .CLK(clk), 
        .QN(n1933) );
  SDFFX1_RVT opC20_d3_reg_12_ ( .D(n3401), .SI(1'b0), .SE(n1982), .CLK(clk), 
        .QN(n1931) );
  SDFFX1_RVT opC20_d3_reg_11_ ( .D(n3401), .SI(1'b0), .SE(n1981), .CLK(clk), 
        .QN(n1929) );
  SDFFX1_RVT opC20_d3_reg_10_ ( .D(n3401), .SI(1'b0), .SE(n1980), .CLK(clk), 
        .QN(n1927) );
  SDFFX1_RVT opC20_d3_reg_9_ ( .D(n3401), .SI(1'b0), .SE(n1979), .CLK(clk), 
        .QN(n1925) );
  SDFFX1_RVT opC20_d3_reg_8_ ( .D(n3401), .SI(1'b0), .SE(n1978), .CLK(clk), 
        .QN(n1923) );
  SDFFX1_RVT opC20_d3_reg_7_ ( .D(n3401), .SI(1'b0), .SE(n1977), .CLK(clk), 
        .QN(n1921) );
  SDFFX1_RVT opC20_d3_reg_6_ ( .D(n3400), .SI(1'b0), .SE(n1976), .CLK(clk), 
        .QN(n1919) );
  SDFFX1_RVT opC20_d3_reg_5_ ( .D(n3400), .SI(1'b0), .SE(n1975), .CLK(clk), 
        .QN(n1917) );
  SDFFX1_RVT opC20_d3_reg_4_ ( .D(n3400), .SI(1'b0), .SE(n1974), .CLK(clk), 
        .QN(n1915) );
  SDFFX1_RVT opC20_d3_reg_3_ ( .D(n3400), .SI(1'b0), .SE(n1973), .CLK(clk), 
        .QN(n1913) );
  SDFFX1_RVT opC20_d3_reg_2_ ( .D(n3400), .SI(1'b0), .SE(n1972), .CLK(clk), 
        .QN(n1911) );
  SDFFX1_RVT opC20_d3_reg_1_ ( .D(n3400), .SI(1'b0), .SE(n1971), .CLK(clk), 
        .QN(n1909) );
  SDFFX1_RVT opC20_d3_reg_0_ ( .D(n3400), .SI(1'b0), .SE(n1970), .CLK(clk), 
        .QN(n1907) );
  SDFFX1_RVT opC20_d2_reg_31_ ( .D(n3400), .SI(1'b0), .SE(n1969), .CLK(clk), 
        .QN(n1905) );
  SDFFX1_RVT opC20_d2_reg_30_ ( .D(n3400), .SI(1'b0), .SE(n1967), .CLK(clk), 
        .QN(n1903) );
  SDFFX1_RVT opC20_d2_reg_29_ ( .D(n3400), .SI(1'b0), .SE(n1965), .CLK(clk), 
        .QN(n1901) );
  SDFFX1_RVT opC20_d2_reg_28_ ( .D(n3400), .SI(1'b0), .SE(n1963), .CLK(clk), 
        .QN(n1899) );
  SDFFX1_RVT opC20_d2_reg_27_ ( .D(n3400), .SI(1'b0), .SE(n1961), .CLK(clk), 
        .QN(n1897) );
  SDFFX1_RVT opC20_d2_reg_26_ ( .D(n3400), .SI(1'b0), .SE(n1959), .CLK(clk), 
        .QN(n1895) );
  SDFFX1_RVT opC20_d2_reg_25_ ( .D(n3400), .SI(1'b0), .SE(n1957), .CLK(clk), 
        .QN(n1893) );
  SDFFX1_RVT opC20_d2_reg_24_ ( .D(n3399), .SI(1'b0), .SE(n1955), .CLK(clk), 
        .QN(n1891) );
  SDFFX1_RVT opC20_d2_reg_23_ ( .D(n3399), .SI(1'b0), .SE(n1953), .CLK(clk), 
        .QN(n1889) );
  SDFFX1_RVT opC20_d2_reg_22_ ( .D(n3399), .SI(1'b0), .SE(n1951), .CLK(clk), 
        .QN(n1887) );
  SDFFX1_RVT opC20_d2_reg_21_ ( .D(n3399), .SI(1'b0), .SE(n1949), .CLK(clk), 
        .QN(n1885) );
  SDFFX1_RVT opC20_d2_reg_20_ ( .D(n3399), .SI(1'b0), .SE(n1947), .CLK(clk), 
        .QN(n1883) );
  SDFFX1_RVT opC20_d2_reg_19_ ( .D(n3399), .SI(1'b0), .SE(n1945), .CLK(clk), 
        .QN(n1881) );
  SDFFX1_RVT opC20_d2_reg_18_ ( .D(n3399), .SI(1'b0), .SE(n1943), .CLK(clk), 
        .QN(n1879) );
  SDFFX1_RVT opC20_d2_reg_17_ ( .D(n3399), .SI(1'b0), .SE(n1941), .CLK(clk), 
        .QN(n1877) );
  SDFFX1_RVT opC20_d2_reg_16_ ( .D(n3399), .SI(1'b0), .SE(n1939), .CLK(clk), 
        .QN(n1875) );
  SDFFX1_RVT opC20_d2_reg_15_ ( .D(n3399), .SI(1'b0), .SE(n1937), .CLK(clk), 
        .QN(n1873) );
  SDFFX1_RVT opC20_d2_reg_14_ ( .D(n3399), .SI(1'b0), .SE(n1935), .CLK(clk), 
        .QN(n1871) );
  SDFFX1_RVT opC20_d2_reg_13_ ( .D(n3403), .SI(1'b0), .SE(n1933), .CLK(clk), 
        .QN(n1869) );
  SDFFX1_RVT opC20_d2_reg_12_ ( .D(n3403), .SI(1'b0), .SE(n1931), .CLK(clk), 
        .QN(n1867) );
  SDFFX1_RVT opC20_d2_reg_11_ ( .D(n3399), .SI(1'b0), .SE(n1929), .CLK(clk), 
        .QN(n1865) );
  SDFFX1_RVT opC20_d2_reg_10_ ( .D(n3399), .SI(1'b0), .SE(n1927), .CLK(clk), 
        .QN(n1863) );
  SDFFX1_RVT opC20_d2_reg_9_ ( .D(n3399), .SI(1'b0), .SE(n1925), .CLK(clk), 
        .QN(n1861) );
  SDFFX1_RVT opC20_d2_reg_8_ ( .D(n3398), .SI(1'b0), .SE(n1923), .CLK(clk), 
        .QN(n1859) );
  SDFFX1_RVT opC20_d2_reg_7_ ( .D(n3398), .SI(1'b0), .SE(n1921), .CLK(clk), 
        .QN(n1857) );
  SDFFX1_RVT opC20_d2_reg_6_ ( .D(n3398), .SI(1'b0), .SE(n1919), .CLK(clk), 
        .QN(n1855) );
  SDFFX1_RVT opC20_d2_reg_5_ ( .D(n3398), .SI(1'b0), .SE(n1917), .CLK(clk), 
        .QN(n1853) );
  SDFFX1_RVT opC20_d2_reg_4_ ( .D(n3398), .SI(1'b0), .SE(n1915), .CLK(clk), 
        .QN(n1851) );
  SDFFX1_RVT opC20_d2_reg_3_ ( .D(n3398), .SI(1'b0), .SE(n1913), .CLK(clk), 
        .QN(n1849) );
  SDFFX1_RVT opC20_d2_reg_2_ ( .D(n3398), .SI(1'b0), .SE(n1911), .CLK(clk), 
        .QN(n1847) );
  SDFFX1_RVT opC20_d2_reg_1_ ( .D(n3398), .SI(1'b0), .SE(n1909), .CLK(clk), 
        .QN(n1845) );
  SDFFX1_RVT opC20_d2_reg_0_ ( .D(n3398), .SI(1'b0), .SE(n1907), .CLK(clk), 
        .QN(n1843) );
  SDFFX1_RVT opC20_d1_reg_31_ ( .D(n3398), .SI(1'b0), .SE(n1905), .CLK(clk), 
        .Q(OpC20[31]) );
  SDFFX1_RVT opC20_d1_reg_30_ ( .D(n3398), .SI(1'b0), .SE(n1903), .CLK(clk), 
        .Q(OpC20[30]) );
  SDFFX1_RVT opC20_d1_reg_29_ ( .D(n3398), .SI(1'b0), .SE(n1901), .CLK(clk), 
        .Q(OpC20[29]) );
  SDFFX1_RVT opC20_d1_reg_28_ ( .D(n3398), .SI(1'b0), .SE(n1899), .CLK(clk), 
        .Q(OpC20[28]) );
  SDFFX1_RVT opC20_d1_reg_27_ ( .D(n3398), .SI(1'b0), .SE(n1897), .CLK(clk), 
        .Q(OpC20[27]) );
  SDFFX1_RVT opC20_d1_reg_26_ ( .D(n3397), .SI(1'b0), .SE(n1895), .CLK(clk), 
        .Q(OpC20[26]) );
  SDFFX1_RVT opC20_d1_reg_25_ ( .D(n3397), .SI(1'b0), .SE(n1893), .CLK(clk), 
        .Q(OpC20[25]) );
  SDFFX1_RVT opC20_d1_reg_24_ ( .D(n3397), .SI(1'b0), .SE(n1891), .CLK(clk), 
        .Q(OpC20[24]) );
  SDFFX1_RVT opC20_d1_reg_23_ ( .D(n3397), .SI(1'b0), .SE(n1889), .CLK(clk), 
        .Q(OpC20[23]) );
  SDFFX1_RVT opC20_d1_reg_22_ ( .D(n3397), .SI(1'b0), .SE(n1887), .CLK(clk), 
        .Q(OpC20[22]) );
  SDFFX1_RVT opC20_d1_reg_21_ ( .D(n3397), .SI(1'b0), .SE(n1885), .CLK(clk), 
        .Q(OpC20[21]) );
  SDFFX1_RVT opC20_d1_reg_20_ ( .D(n3397), .SI(1'b0), .SE(n1883), .CLK(clk), 
        .Q(OpC20[20]) );
  SDFFX1_RVT opC20_d1_reg_19_ ( .D(n3397), .SI(1'b0), .SE(n1881), .CLK(clk), 
        .Q(OpC20[19]) );
  SDFFX1_RVT opC20_d1_reg_18_ ( .D(n3397), .SI(1'b0), .SE(n1879), .CLK(clk), 
        .Q(OpC20[18]) );
  SDFFX1_RVT opC20_d1_reg_17_ ( .D(n3397), .SI(1'b0), .SE(n1877), .CLK(clk), 
        .Q(OpC20[17]) );
  SDFFX1_RVT opC20_d1_reg_16_ ( .D(n3397), .SI(1'b0), .SE(n1875), .CLK(clk), 
        .Q(OpC20[16]) );
  SDFFX1_RVT opC20_d1_reg_15_ ( .D(n3397), .SI(1'b0), .SE(n1873), .CLK(clk), 
        .Q(OpC20[15]) );
  SDFFX1_RVT opC20_d1_reg_14_ ( .D(n3397), .SI(1'b0), .SE(n1871), .CLK(clk), 
        .Q(OpC20[14]) );
  SDFFX1_RVT opC20_d1_reg_13_ ( .D(n3397), .SI(1'b0), .SE(n1869), .CLK(clk), 
        .Q(OpC20[13]) );
  SDFFX1_RVT opC20_d1_reg_12_ ( .D(n3396), .SI(1'b0), .SE(n1867), .CLK(clk), 
        .Q(OpC20[12]) );
  SDFFX1_RVT opC20_d1_reg_11_ ( .D(n3396), .SI(1'b0), .SE(n1865), .CLK(clk), 
        .Q(OpC20[11]) );
  SDFFX1_RVT opC20_d1_reg_10_ ( .D(n3396), .SI(1'b0), .SE(n1863), .CLK(clk), 
        .Q(OpC20[10]) );
  SDFFX1_RVT opC20_d1_reg_9_ ( .D(n3396), .SI(1'b0), .SE(n1861), .CLK(clk), 
        .Q(OpC20[9]) );
  SDFFX1_RVT opC20_d1_reg_8_ ( .D(n3396), .SI(1'b0), .SE(n1859), .CLK(clk), 
        .Q(OpC20[8]) );
  SDFFX1_RVT opC20_d1_reg_7_ ( .D(n3396), .SI(1'b0), .SE(n1857), .CLK(clk), 
        .Q(OpC20[7]) );
  SDFFX1_RVT opC20_d1_reg_6_ ( .D(n3396), .SI(1'b0), .SE(n1855), .CLK(clk), 
        .Q(OpC20[6]) );
  SDFFX1_RVT opC20_d1_reg_5_ ( .D(n3396), .SI(1'b0), .SE(n1853), .CLK(clk), 
        .Q(OpC20[5]) );
  SDFFX1_RVT opC20_d1_reg_4_ ( .D(n3396), .SI(1'b0), .SE(n1851), .CLK(clk), 
        .Q(OpC20[4]) );
  SDFFX1_RVT opC20_d1_reg_3_ ( .D(n3396), .SI(1'b0), .SE(n1849), .CLK(clk), 
        .Q(OpC20[3]) );
  SDFFX1_RVT opC20_d1_reg_2_ ( .D(n3396), .SI(1'b0), .SE(n1847), .CLK(clk), 
        .Q(OpC20[2]) );
  SDFFX1_RVT opC20_d1_reg_1_ ( .D(n3396), .SI(1'b0), .SE(n1845), .CLK(clk), 
        .Q(OpC20[1]) );
  SDFFX1_RVT opC20_d1_reg_0_ ( .D(n3396), .SI(1'b0), .SE(n1843), .CLK(clk), 
        .Q(OpC20[0]) );
  SDFFX1_RVT opC03_d2_reg_31_ ( .D(n3396), .SI(1'b0), .SE(n1809), .CLK(clk), 
        .QN(n1777) );
  SDFFX1_RVT opC03_d2_reg_30_ ( .D(n3395), .SI(1'b0), .SE(n1808), .CLK(clk), 
        .QN(n1775) );
  SDFFX1_RVT opC03_d2_reg_29_ ( .D(n3395), .SI(1'b0), .SE(n1807), .CLK(clk), 
        .QN(n1773) );
  SDFFX1_RVT opC03_d2_reg_28_ ( .D(n3395), .SI(1'b0), .SE(n1806), .CLK(clk), 
        .QN(n1771) );
  SDFFX1_RVT opC03_d2_reg_27_ ( .D(n3395), .SI(1'b0), .SE(n1805), .CLK(clk), 
        .QN(n1769) );
  SDFFX1_RVT opC03_d2_reg_26_ ( .D(n3395), .SI(1'b0), .SE(n1804), .CLK(clk), 
        .QN(n1767) );
  SDFFX1_RVT opC03_d2_reg_25_ ( .D(n3395), .SI(1'b0), .SE(n1803), .CLK(clk), 
        .QN(n1765) );
  SDFFX1_RVT opC03_d2_reg_24_ ( .D(n3395), .SI(1'b0), .SE(n1802), .CLK(clk), 
        .QN(n1763) );
  SDFFX1_RVT opC03_d2_reg_23_ ( .D(n3395), .SI(1'b0), .SE(n1801), .CLK(clk), 
        .QN(n1761) );
  SDFFX1_RVT opC03_d2_reg_22_ ( .D(n3395), .SI(1'b0), .SE(n1800), .CLK(clk), 
        .QN(n1759) );
  SDFFX1_RVT opC03_d2_reg_21_ ( .D(n3395), .SI(1'b0), .SE(n1799), .CLK(clk), 
        .QN(n1757) );
  SDFFX1_RVT opC03_d2_reg_20_ ( .D(n3395), .SI(1'b0), .SE(n1798), .CLK(clk), 
        .QN(n1755) );
  SDFFX1_RVT opC03_d2_reg_19_ ( .D(n3395), .SI(1'b0), .SE(n1797), .CLK(clk), 
        .QN(n1753) );
  SDFFX1_RVT opC03_d2_reg_18_ ( .D(n3395), .SI(1'b0), .SE(n1796), .CLK(clk), 
        .QN(n1751) );
  SDFFX1_RVT opC03_d2_reg_17_ ( .D(n3395), .SI(1'b0), .SE(n1795), .CLK(clk), 
        .QN(n1749) );
  SDFFX1_RVT opC03_d2_reg_16_ ( .D(n3394), .SI(1'b0), .SE(n1794), .CLK(clk), 
        .QN(n1747) );
  SDFFX1_RVT opC03_d2_reg_15_ ( .D(n3394), .SI(1'b0), .SE(n1793), .CLK(clk), 
        .QN(n1745) );
  SDFFX1_RVT opC03_d2_reg_14_ ( .D(n3394), .SI(1'b0), .SE(n1792), .CLK(clk), 
        .QN(n1743) );
  SDFFX1_RVT opC03_d2_reg_13_ ( .D(n3394), .SI(1'b0), .SE(n1791), .CLK(clk), 
        .QN(n1741) );
  SDFFX1_RVT opC03_d2_reg_12_ ( .D(n3394), .SI(1'b0), .SE(n1790), .CLK(clk), 
        .QN(n1739) );
  SDFFX1_RVT opC03_d2_reg_11_ ( .D(n3394), .SI(1'b0), .SE(n1789), .CLK(clk), 
        .QN(n1737) );
  SDFFX1_RVT opC03_d2_reg_10_ ( .D(n3394), .SI(1'b0), .SE(n1788), .CLK(clk), 
        .QN(n1735) );
  SDFFX1_RVT opC03_d2_reg_9_ ( .D(n3394), .SI(1'b0), .SE(n1787), .CLK(clk), 
        .QN(n1733) );
  SDFFX1_RVT opC03_d2_reg_8_ ( .D(n3394), .SI(1'b0), .SE(n1786), .CLK(clk), 
        .QN(n1731) );
  SDFFX1_RVT opC03_d2_reg_7_ ( .D(n3394), .SI(1'b0), .SE(n1785), .CLK(clk), 
        .QN(n1729) );
  SDFFX1_RVT opC03_d2_reg_6_ ( .D(n3394), .SI(1'b0), .SE(n1784), .CLK(clk), 
        .QN(n1727) );
  SDFFX1_RVT opC03_d2_reg_5_ ( .D(n3394), .SI(1'b0), .SE(n1783), .CLK(clk), 
        .QN(n1725) );
  SDFFX1_RVT opC03_d2_reg_4_ ( .D(n3393), .SI(1'b0), .SE(n1782), .CLK(clk), 
        .QN(n1723) );
  SDFFX1_RVT opC03_d2_reg_3_ ( .D(n3393), .SI(1'b0), .SE(n1781), .CLK(clk), 
        .QN(n1721) );
  SDFFX1_RVT opC03_d2_reg_2_ ( .D(n3393), .SI(1'b0), .SE(n1780), .CLK(clk), 
        .QN(n1719) );
  SDFFX1_RVT opC03_d2_reg_1_ ( .D(n3393), .SI(1'b0), .SE(n1779), .CLK(clk), 
        .QN(n1717) );
  SDFFX1_RVT opC03_d2_reg_0_ ( .D(n3393), .SI(1'b0), .SE(n1778), .CLK(clk), 
        .QN(n1715) );
  SDFFX1_RVT opC03_d1_reg_31_ ( .D(n3393), .SI(1'b0), .SE(n1777), .CLK(clk), 
        .Q(OpC03[31]) );
  SDFFX1_RVT opC03_d1_reg_30_ ( .D(n3393), .SI(1'b0), .SE(n1775), .CLK(clk), 
        .Q(OpC03[30]) );
  SDFFX1_RVT opC03_d1_reg_29_ ( .D(n3393), .SI(1'b0), .SE(n1773), .CLK(clk), 
        .Q(OpC03[29]) );
  SDFFX1_RVT opC03_d1_reg_28_ ( .D(n3393), .SI(1'b0), .SE(n1771), .CLK(clk), 
        .Q(OpC03[28]) );
  SDFFX1_RVT opC03_d1_reg_27_ ( .D(n3393), .SI(1'b0), .SE(n1769), .CLK(clk), 
        .Q(OpC03[27]) );
  SDFFX1_RVT opC03_d1_reg_26_ ( .D(n3393), .SI(1'b0), .SE(n1767), .CLK(clk), 
        .Q(OpC03[26]) );
  SDFFX1_RVT opC03_d1_reg_25_ ( .D(n3393), .SI(1'b0), .SE(n1765), .CLK(clk), 
        .Q(OpC03[25]) );
  SDFFX1_RVT opC03_d1_reg_24_ ( .D(n3393), .SI(1'b0), .SE(n1763), .CLK(clk), 
        .Q(OpC03[24]) );
  SDFFX1_RVT opC03_d1_reg_23_ ( .D(n3393), .SI(1'b0), .SE(n1761), .CLK(clk), 
        .Q(OpC03[23]) );
  SDFFX1_RVT opC03_d1_reg_22_ ( .D(n3392), .SI(1'b0), .SE(n1759), .CLK(clk), 
        .Q(OpC03[22]) );
  SDFFX1_RVT opC03_d1_reg_21_ ( .D(n3392), .SI(1'b0), .SE(n1757), .CLK(clk), 
        .Q(OpC03[21]) );
  SDFFX1_RVT opC03_d1_reg_20_ ( .D(n3392), .SI(1'b0), .SE(n1755), .CLK(clk), 
        .Q(OpC03[20]) );
  SDFFX1_RVT opC03_d1_reg_19_ ( .D(n3392), .SI(1'b0), .SE(n1753), .CLK(clk), 
        .Q(OpC03[19]) );
  SDFFX1_RVT opC03_d1_reg_18_ ( .D(n3392), .SI(1'b0), .SE(n1751), .CLK(clk), 
        .Q(OpC03[18]) );
  SDFFX1_RVT opC03_d1_reg_17_ ( .D(n3392), .SI(1'b0), .SE(n1749), .CLK(clk), 
        .Q(OpC03[17]) );
  SDFFX1_RVT opC03_d1_reg_16_ ( .D(n3392), .SI(1'b0), .SE(n1747), .CLK(clk), 
        .Q(OpC03[16]) );
  SDFFX1_RVT opC03_d1_reg_15_ ( .D(n3392), .SI(1'b0), .SE(n1745), .CLK(clk), 
        .Q(OpC03[15]) );
  SDFFX1_RVT opC03_d1_reg_14_ ( .D(n3392), .SI(1'b0), .SE(n1743), .CLK(clk), 
        .Q(OpC03[14]) );
  SDFFX1_RVT opC03_d1_reg_13_ ( .D(n3392), .SI(1'b0), .SE(n1741), .CLK(clk), 
        .Q(OpC03[13]) );
  SDFFX1_RVT opC03_d1_reg_12_ ( .D(n3392), .SI(1'b0), .SE(n1739), .CLK(clk), 
        .Q(OpC03[12]) );
  SDFFX1_RVT opC03_d1_reg_11_ ( .D(n3392), .SI(1'b0), .SE(n1737), .CLK(clk), 
        .Q(OpC03[11]) );
  SDFFX1_RVT opC03_d1_reg_10_ ( .D(n3392), .SI(1'b0), .SE(n1735), .CLK(clk), 
        .Q(OpC03[10]) );
  SDFFX1_RVT opC03_d1_reg_9_ ( .D(n3392), .SI(1'b0), .SE(n1733), .CLK(clk), 
        .Q(OpC03[9]) );
  SDFFX1_RVT opC03_d1_reg_8_ ( .D(n3391), .SI(1'b0), .SE(n1731), .CLK(clk), 
        .Q(OpC03[8]) );
  SDFFX1_RVT opC03_d1_reg_7_ ( .D(n3391), .SI(1'b0), .SE(n1729), .CLK(clk), 
        .Q(OpC03[7]) );
  SDFFX1_RVT opC03_d1_reg_6_ ( .D(n3391), .SI(1'b0), .SE(n1727), .CLK(clk), 
        .Q(OpC03[6]) );
  SDFFX1_RVT opC03_d1_reg_5_ ( .D(n3391), .SI(1'b0), .SE(n1725), .CLK(clk), 
        .Q(OpC03[5]) );
  SDFFX1_RVT opC03_d1_reg_4_ ( .D(n3391), .SI(1'b0), .SE(n1723), .CLK(clk), 
        .Q(OpC03[4]) );
  SDFFX1_RVT opC03_d1_reg_3_ ( .D(n3391), .SI(1'b0), .SE(n1721), .CLK(clk), 
        .Q(OpC03[3]) );
  SDFFX1_RVT opC03_d1_reg_2_ ( .D(n3391), .SI(1'b0), .SE(n1719), .CLK(clk), 
        .Q(OpC03[2]) );
  SDFFX1_RVT opC03_d1_reg_1_ ( .D(n3391), .SI(1'b0), .SE(n1717), .CLK(clk), 
        .Q(OpC03[1]) );
  SDFFX1_RVT opC03_d1_reg_0_ ( .D(n3391), .SI(1'b0), .SE(n1715), .CLK(clk), 
        .Q(OpC03[0]) );
  SDFFX1_RVT opC12_d2_reg_31_ ( .D(n3391), .SI(1'b0), .SE(n1681), .CLK(clk), 
        .QN(n1649) );
  SDFFX1_RVT opC12_d2_reg_30_ ( .D(n3391), .SI(1'b0), .SE(n1680), .CLK(clk), 
        .QN(n1647) );
  SDFFX1_RVT opC12_d2_reg_29_ ( .D(n3391), .SI(1'b0), .SE(n1679), .CLK(clk), 
        .QN(n1645) );
  SDFFX1_RVT opC12_d2_reg_28_ ( .D(n3391), .SI(1'b0), .SE(n1678), .CLK(clk), 
        .QN(n1643) );
  SDFFX1_RVT opC12_d2_reg_27_ ( .D(n3391), .SI(1'b0), .SE(n1677), .CLK(clk), 
        .QN(n1641) );
  SDFFX1_RVT opC12_d2_reg_26_ ( .D(n3475), .SI(1'b0), .SE(n1676), .CLK(clk), 
        .QN(n1639) );
  SDFFX1_RVT opC12_d2_reg_25_ ( .D(n3474), .SI(1'b0), .SE(n1675), .CLK(clk), 
        .QN(n1637) );
  SDFFX1_RVT opC12_d2_reg_24_ ( .D(n3475), .SI(1'b0), .SE(n1674), .CLK(clk), 
        .QN(n1635) );
  SDFFX1_RVT opC12_d2_reg_23_ ( .D(n3474), .SI(1'b0), .SE(n1673), .CLK(clk), 
        .QN(n1633) );
  SDFFX1_RVT opC12_d2_reg_22_ ( .D(n3475), .SI(1'b0), .SE(n1672), .CLK(clk), 
        .QN(n1631) );
  SDFFX1_RVT opC12_d2_reg_21_ ( .D(n3474), .SI(1'b0), .SE(n1671), .CLK(clk), 
        .QN(n1629) );
  SDFFX1_RVT opC12_d2_reg_20_ ( .D(n3475), .SI(1'b0), .SE(n1670), .CLK(clk), 
        .QN(n1627) );
  SDFFX1_RVT opC12_d2_reg_19_ ( .D(n3462), .SI(1'b0), .SE(n1669), .CLK(clk), 
        .QN(n1625) );
  SDFFX1_RVT opC12_d2_reg_18_ ( .D(n3461), .SI(1'b0), .SE(n1668), .CLK(clk), 
        .QN(n1623) );
  SDFFX1_RVT opC12_d2_reg_17_ ( .D(n3463), .SI(1'b0), .SE(n1667), .CLK(clk), 
        .QN(n1621) );
  SDFFX1_RVT opC12_d2_reg_16_ ( .D(n3459), .SI(1'b0), .SE(n1666), .CLK(clk), 
        .QN(n1619) );
  SDFFX1_RVT opC12_d2_reg_15_ ( .D(n3460), .SI(1'b0), .SE(n1665), .CLK(clk), 
        .QN(n1617) );
  SDFFX1_RVT opC12_d2_reg_14_ ( .D(n3458), .SI(1'b0), .SE(n1664), .CLK(clk), 
        .QN(n1615) );
  SDFFX1_RVT opC12_d2_reg_13_ ( .D(n3458), .SI(1'b0), .SE(n1663), .CLK(clk), 
        .QN(n1613) );
  SDFFX1_RVT opC12_d2_reg_12_ ( .D(n3390), .SI(1'b0), .SE(n1662), .CLK(clk), 
        .QN(n1611) );
  SDFFX1_RVT opC12_d2_reg_11_ ( .D(n3390), .SI(1'b0), .SE(n1661), .CLK(clk), 
        .QN(n1609) );
  SDFFX1_RVT opC12_d2_reg_10_ ( .D(n3390), .SI(1'b0), .SE(n1660), .CLK(clk), 
        .QN(n1607) );
  SDFFX1_RVT opC12_d2_reg_9_ ( .D(n3394), .SI(1'b0), .SE(n1659), .CLK(clk), 
        .QN(n1605) );
  SDFFX1_RVT opC12_d2_reg_8_ ( .D(n3390), .SI(1'b0), .SE(n1658), .CLK(clk), 
        .QN(n1603) );
  SDFFX1_RVT opC12_d2_reg_7_ ( .D(n3390), .SI(1'b0), .SE(n1657), .CLK(clk), 
        .QN(n1601) );
  SDFFX1_RVT opC12_d2_reg_6_ ( .D(n3390), .SI(1'b0), .SE(n1656), .CLK(clk), 
        .QN(n1599) );
  SDFFX1_RVT opC12_d2_reg_5_ ( .D(n3390), .SI(1'b0), .SE(n1655), .CLK(clk), 
        .QN(n1597) );
  SDFFX1_RVT opC12_d2_reg_4_ ( .D(n3390), .SI(1'b0), .SE(n1654), .CLK(clk), 
        .QN(n1595) );
  SDFFX1_RVT opC12_d2_reg_3_ ( .D(n3390), .SI(1'b0), .SE(n1653), .CLK(clk), 
        .QN(n1593) );
  SDFFX1_RVT opC12_d2_reg_2_ ( .D(n3390), .SI(1'b0), .SE(n1652), .CLK(clk), 
        .QN(n1591) );
  SDFFX1_RVT opC12_d2_reg_1_ ( .D(n3390), .SI(1'b0), .SE(n1651), .CLK(clk), 
        .QN(n1589) );
  SDFFX1_RVT opC12_d2_reg_0_ ( .D(n3390), .SI(1'b0), .SE(n1650), .CLK(clk), 
        .QN(n1587) );
  SDFFX1_RVT opC12_d1_reg_31_ ( .D(n3390), .SI(1'b0), .SE(n1649), .CLK(clk), 
        .Q(OpC12[31]) );
  SDFFX1_RVT opC12_d1_reg_30_ ( .D(n3389), .SI(1'b0), .SE(n1647), .CLK(clk), 
        .Q(OpC12[30]) );
  SDFFX1_RVT opC12_d1_reg_29_ ( .D(n3389), .SI(1'b0), .SE(n1645), .CLK(clk), 
        .Q(OpC12[29]) );
  SDFFX1_RVT opC12_d1_reg_28_ ( .D(n3389), .SI(1'b0), .SE(n1643), .CLK(clk), 
        .Q(OpC12[28]) );
  SDFFX1_RVT opC12_d1_reg_27_ ( .D(n3389), .SI(1'b0), .SE(n1641), .CLK(clk), 
        .Q(OpC12[27]) );
  SDFFX1_RVT opC12_d1_reg_26_ ( .D(n3389), .SI(1'b0), .SE(n1639), .CLK(clk), 
        .Q(OpC12[26]) );
  SDFFX1_RVT opC12_d1_reg_25_ ( .D(n3389), .SI(1'b0), .SE(n1637), .CLK(clk), 
        .Q(OpC12[25]) );
  SDFFX1_RVT opC12_d1_reg_24_ ( .D(n3389), .SI(1'b0), .SE(n1635), .CLK(clk), 
        .Q(OpC12[24]) );
  SDFFX1_RVT opC12_d1_reg_23_ ( .D(n3389), .SI(1'b0), .SE(n1633), .CLK(clk), 
        .Q(OpC12[23]) );
  SDFFX1_RVT opC12_d1_reg_22_ ( .D(n3389), .SI(1'b0), .SE(n1631), .CLK(clk), 
        .Q(OpC12[22]) );
  SDFFX1_RVT opC12_d1_reg_21_ ( .D(n3389), .SI(1'b0), .SE(n1629), .CLK(clk), 
        .Q(OpC12[21]) );
  SDFFX1_RVT opC12_d1_reg_20_ ( .D(n3389), .SI(1'b0), .SE(n1627), .CLK(clk), 
        .Q(OpC12[20]) );
  SDFFX1_RVT opC12_d1_reg_19_ ( .D(n3389), .SI(1'b0), .SE(n1625), .CLK(clk), 
        .Q(OpC12[19]) );
  SDFFX1_RVT opC12_d1_reg_18_ ( .D(n3389), .SI(1'b0), .SE(n1623), .CLK(clk), 
        .Q(OpC12[18]) );
  SDFFX1_RVT opC12_d1_reg_17_ ( .D(n3389), .SI(1'b0), .SE(n1621), .CLK(clk), 
        .Q(OpC12[17]) );
  SDFFX1_RVT opC12_d1_reg_16_ ( .D(n3388), .SI(1'b0), .SE(n1619), .CLK(clk), 
        .Q(OpC12[16]) );
  SDFFX1_RVT opC12_d1_reg_15_ ( .D(n3388), .SI(1'b0), .SE(n1617), .CLK(clk), 
        .Q(OpC12[15]) );
  SDFFX1_RVT opC12_d1_reg_14_ ( .D(n3388), .SI(1'b0), .SE(n1615), .CLK(clk), 
        .Q(OpC12[14]) );
  SDFFX1_RVT opC12_d1_reg_13_ ( .D(n3388), .SI(1'b0), .SE(n1613), .CLK(clk), 
        .Q(OpC12[13]) );
  SDFFX1_RVT opC12_d1_reg_12_ ( .D(n3388), .SI(1'b0), .SE(n1611), .CLK(clk), 
        .Q(OpC12[12]) );
  SDFFX1_RVT opC12_d1_reg_11_ ( .D(n3388), .SI(1'b0), .SE(n1609), .CLK(clk), 
        .Q(OpC12[11]) );
  SDFFX1_RVT opC12_d1_reg_10_ ( .D(n3388), .SI(1'b0), .SE(n1607), .CLK(clk), 
        .Q(OpC12[10]) );
  SDFFX1_RVT opC12_d1_reg_9_ ( .D(n3388), .SI(1'b0), .SE(n1605), .CLK(clk), 
        .Q(OpC12[9]) );
  SDFFX1_RVT opC12_d1_reg_8_ ( .D(n3388), .SI(1'b0), .SE(n1603), .CLK(clk), 
        .Q(OpC12[8]) );
  SDFFX1_RVT opC12_d1_reg_7_ ( .D(n3388), .SI(1'b0), .SE(n1601), .CLK(clk), 
        .Q(OpC12[7]) );
  SDFFX1_RVT opC12_d1_reg_6_ ( .D(n3388), .SI(1'b0), .SE(n1599), .CLK(clk), 
        .Q(OpC12[6]) );
  SDFFX1_RVT opC12_d1_reg_5_ ( .D(n3388), .SI(1'b0), .SE(n1597), .CLK(clk), 
        .Q(OpC12[5]) );
  SDFFX1_RVT opC12_d1_reg_4_ ( .D(n3388), .SI(1'b0), .SE(n1595), .CLK(clk), 
        .Q(OpC12[4]) );
  SDFFX1_RVT opC12_d1_reg_3_ ( .D(n3388), .SI(1'b0), .SE(n1593), .CLK(clk), 
        .Q(OpC12[3]) );
  SDFFX1_RVT opC12_d1_reg_2_ ( .D(n3387), .SI(1'b0), .SE(n1591), .CLK(clk), 
        .Q(OpC12[2]) );
  SDFFX1_RVT opC12_d1_reg_1_ ( .D(n3387), .SI(1'b0), .SE(n1589), .CLK(clk), 
        .Q(OpC12[1]) );
  SDFFX1_RVT opC12_d1_reg_0_ ( .D(n3387), .SI(1'b0), .SE(n1587), .CLK(clk), 
        .Q(OpC12[0]) );
  SDFFX1_RVT opC21_d2_reg_31_ ( .D(n3387), .SI(1'b0), .SE(n1553), .CLK(clk), 
        .QN(n1521) );
  SDFFX1_RVT opC21_d2_reg_30_ ( .D(n3387), .SI(1'b0), .SE(n1552), .CLK(clk), 
        .QN(n1519) );
  SDFFX1_RVT opC21_d2_reg_29_ ( .D(n3387), .SI(1'b0), .SE(n1551), .CLK(clk), 
        .QN(n1517) );
  SDFFX1_RVT opC21_d2_reg_28_ ( .D(n3387), .SI(1'b0), .SE(n1550), .CLK(clk), 
        .QN(n1515) );
  SDFFX1_RVT opC21_d2_reg_27_ ( .D(n3387), .SI(1'b0), .SE(n1549), .CLK(clk), 
        .QN(n1513) );
  SDFFX1_RVT opC21_d2_reg_26_ ( .D(n3387), .SI(1'b0), .SE(n1548), .CLK(clk), 
        .QN(n1511) );
  SDFFX1_RVT opC21_d2_reg_25_ ( .D(n3387), .SI(1'b0), .SE(n1547), .CLK(clk), 
        .QN(n1509) );
  SDFFX1_RVT opC21_d2_reg_24_ ( .D(n3387), .SI(1'b0), .SE(n1546), .CLK(clk), 
        .QN(n1507) );
  SDFFX1_RVT opC21_d2_reg_23_ ( .D(n3387), .SI(1'b0), .SE(n1545), .CLK(clk), 
        .QN(n1505) );
  SDFFX1_RVT opC21_d2_reg_22_ ( .D(n3387), .SI(1'b0), .SE(n1544), .CLK(clk), 
        .QN(n1503) );
  SDFFX1_RVT opC21_d2_reg_21_ ( .D(n3387), .SI(1'b0), .SE(n1543), .CLK(clk), 
        .QN(n1501) );
  SDFFX1_RVT opC21_d2_reg_20_ ( .D(n3386), .SI(1'b0), .SE(n1542), .CLK(clk), 
        .QN(n1499) );
  SDFFX1_RVT opC21_d2_reg_19_ ( .D(n3386), .SI(1'b0), .SE(n1541), .CLK(clk), 
        .QN(n1497) );
  SDFFX1_RVT opC21_d2_reg_18_ ( .D(n3386), .SI(1'b0), .SE(n1540), .CLK(clk), 
        .QN(n1495) );
  SDFFX1_RVT opC21_d2_reg_17_ ( .D(n3386), .SI(1'b0), .SE(n1539), .CLK(clk), 
        .QN(n1493) );
  SDFFX1_RVT opC21_d2_reg_16_ ( .D(n3386), .SI(1'b0), .SE(n1538), .CLK(clk), 
        .QN(n1491) );
  SDFFX1_RVT opC21_d2_reg_15_ ( .D(n3386), .SI(1'b0), .SE(n1537), .CLK(clk), 
        .QN(n1489) );
  SDFFX1_RVT opC21_d2_reg_14_ ( .D(n3386), .SI(1'b0), .SE(n1536), .CLK(clk), 
        .QN(n1487) );
  SDFFX1_RVT opC21_d2_reg_13_ ( .D(n3386), .SI(1'b0), .SE(n1535), .CLK(clk), 
        .QN(n1485) );
  SDFFX1_RVT opC21_d2_reg_12_ ( .D(n3386), .SI(1'b0), .SE(n1534), .CLK(clk), 
        .QN(n1483) );
  SDFFX1_RVT opC21_d2_reg_11_ ( .D(n3386), .SI(1'b0), .SE(n1533), .CLK(clk), 
        .QN(n1481) );
  SDFFX1_RVT opC21_d2_reg_10_ ( .D(n3386), .SI(1'b0), .SE(n1532), .CLK(clk), 
        .QN(n1479) );
  SDFFX1_RVT opC21_d2_reg_9_ ( .D(n3386), .SI(1'b0), .SE(n1531), .CLK(clk), 
        .QN(n1477) );
  SDFFX1_RVT opC21_d2_reg_8_ ( .D(n3386), .SI(1'b0), .SE(n1530), .CLK(clk), 
        .QN(n1475) );
  SDFFX1_RVT opC21_d2_reg_7_ ( .D(n3385), .SI(1'b0), .SE(n1529), .CLK(clk), 
        .QN(n1473) );
  SDFFX1_RVT opC21_d2_reg_6_ ( .D(n3385), .SI(1'b0), .SE(n1528), .CLK(clk), 
        .QN(n1471) );
  SDFFX1_RVT opC21_d2_reg_5_ ( .D(n3385), .SI(1'b0), .SE(n1527), .CLK(clk), 
        .QN(n1469) );
  SDFFX1_RVT opC21_d2_reg_4_ ( .D(n3385), .SI(1'b0), .SE(n1526), .CLK(clk), 
        .QN(n1467) );
  SDFFX1_RVT opC21_d2_reg_3_ ( .D(n3385), .SI(1'b0), .SE(n1525), .CLK(clk), 
        .QN(n1465) );
  SDFFX1_RVT opC21_d2_reg_2_ ( .D(n3385), .SI(1'b0), .SE(n1524), .CLK(clk), 
        .QN(n1463) );
  SDFFX1_RVT opC21_d2_reg_1_ ( .D(n3385), .SI(1'b0), .SE(n1523), .CLK(clk), 
        .QN(n1461) );
  SDFFX1_RVT opC21_d2_reg_0_ ( .D(n3385), .SI(1'b0), .SE(n1522), .CLK(clk), 
        .QN(n1459) );
  SDFFX1_RVT opC21_d1_reg_31_ ( .D(n3385), .SI(1'b0), .SE(n1521), .CLK(clk), 
        .Q(OpC21[31]) );
  SDFFX1_RVT opC21_d1_reg_30_ ( .D(n3385), .SI(1'b0), .SE(n1519), .CLK(clk), 
        .Q(OpC21[30]) );
  SDFFX1_RVT opC21_d1_reg_29_ ( .D(n3385), .SI(1'b0), .SE(n1517), .CLK(clk), 
        .Q(OpC21[29]) );
  SDFFX1_RVT opC21_d1_reg_28_ ( .D(n3385), .SI(1'b0), .SE(n1515), .CLK(clk), 
        .Q(OpC21[28]) );
  SDFFX1_RVT opC21_d1_reg_27_ ( .D(n3385), .SI(1'b0), .SE(n1513), .CLK(clk), 
        .Q(OpC21[27]) );
  SDFFX1_RVT opC21_d1_reg_26_ ( .D(n3384), .SI(1'b0), .SE(n1511), .CLK(clk), 
        .Q(OpC21[26]) );
  SDFFX1_RVT opC21_d1_reg_25_ ( .D(n3384), .SI(1'b0), .SE(n1509), .CLK(clk), 
        .Q(OpC21[25]) );
  SDFFX1_RVT opC21_d1_reg_24_ ( .D(n3384), .SI(1'b0), .SE(n1507), .CLK(clk), 
        .Q(OpC21[24]) );
  SDFFX1_RVT opC21_d1_reg_23_ ( .D(n3384), .SI(1'b0), .SE(n1505), .CLK(clk), 
        .Q(OpC21[23]) );
  SDFFX1_RVT opC21_d1_reg_22_ ( .D(n3384), .SI(1'b0), .SE(n1503), .CLK(clk), 
        .Q(OpC21[22]) );
  SDFFX1_RVT opC21_d1_reg_21_ ( .D(n3384), .SI(1'b0), .SE(n1501), .CLK(clk), 
        .Q(OpC21[21]) );
  SDFFX1_RVT opC21_d1_reg_20_ ( .D(n3384), .SI(1'b0), .SE(n1499), .CLK(clk), 
        .Q(OpC21[20]) );
  SDFFX1_RVT opC21_d1_reg_19_ ( .D(n3384), .SI(1'b0), .SE(n1497), .CLK(clk), 
        .Q(OpC21[19]) );
  SDFFX1_RVT opC21_d1_reg_18_ ( .D(n3384), .SI(1'b0), .SE(n1495), .CLK(clk), 
        .Q(OpC21[18]) );
  SDFFX1_RVT opC21_d1_reg_17_ ( .D(n3384), .SI(1'b0), .SE(n1493), .CLK(clk), 
        .Q(OpC21[17]) );
  SDFFX1_RVT opC21_d1_reg_16_ ( .D(n3384), .SI(1'b0), .SE(n1491), .CLK(clk), 
        .Q(OpC21[16]) );
  SDFFX1_RVT opC21_d1_reg_15_ ( .D(n3384), .SI(1'b0), .SE(n1489), .CLK(clk), 
        .Q(OpC21[15]) );
  SDFFX1_RVT opC21_d1_reg_14_ ( .D(n3384), .SI(1'b0), .SE(n1487), .CLK(clk), 
        .Q(OpC21[14]) );
  SDFFX1_RVT opC21_d1_reg_13_ ( .D(n3384), .SI(1'b0), .SE(n1485), .CLK(clk), 
        .Q(OpC21[13]) );
  SDFFX1_RVT opC21_d1_reg_12_ ( .D(n3383), .SI(1'b0), .SE(n1483), .CLK(clk), 
        .Q(OpC21[12]) );
  SDFFX1_RVT opC21_d1_reg_11_ ( .D(n3383), .SI(1'b0), .SE(n1481), .CLK(clk), 
        .Q(OpC21[11]) );
  SDFFX1_RVT opC21_d1_reg_10_ ( .D(n3383), .SI(1'b0), .SE(n1479), .CLK(clk), 
        .Q(OpC21[10]) );
  SDFFX1_RVT opC21_d1_reg_9_ ( .D(n3383), .SI(1'b0), .SE(n1477), .CLK(clk), 
        .Q(OpC21[9]) );
  SDFFX1_RVT opC21_d1_reg_8_ ( .D(n3383), .SI(1'b0), .SE(n1475), .CLK(clk), 
        .Q(OpC21[8]) );
  SDFFX1_RVT opC21_d1_reg_7_ ( .D(n3383), .SI(1'b0), .SE(n1473), .CLK(clk), 
        .Q(OpC21[7]) );
  SDFFX1_RVT opC21_d1_reg_6_ ( .D(n3383), .SI(1'b0), .SE(n1471), .CLK(clk), 
        .Q(OpC21[6]) );
  SDFFX1_RVT opC21_d1_reg_5_ ( .D(n3383), .SI(1'b0), .SE(n1469), .CLK(clk), 
        .Q(OpC21[5]) );
  SDFFX1_RVT opC21_d1_reg_4_ ( .D(n3383), .SI(1'b0), .SE(n1467), .CLK(clk), 
        .Q(OpC21[4]) );
  SDFFX1_RVT opC21_d1_reg_3_ ( .D(n3383), .SI(1'b0), .SE(n1465), .CLK(clk), 
        .Q(OpC21[3]) );
  SDFFX1_RVT opC21_d1_reg_2_ ( .D(n3383), .SI(1'b0), .SE(n1463), .CLK(clk), 
        .Q(OpC21[2]) );
  SDFFX1_RVT opC21_d1_reg_1_ ( .D(n3383), .SI(1'b0), .SE(n1461), .CLK(clk), 
        .Q(OpC21[1]) );
  SDFFX1_RVT opC21_d1_reg_0_ ( .D(n3383), .SI(1'b0), .SE(n1459), .CLK(clk), 
        .Q(OpC21[0]) );
  SDFFX1_RVT opC30_d2_reg_31_ ( .D(n3383), .SI(1'b0), .SE(n1425), .CLK(clk), 
        .QN(n1393) );
  SDFFX1_RVT opC30_d2_reg_30_ ( .D(n3382), .SI(1'b0), .SE(n1424), .CLK(clk), 
        .QN(n1391) );
  SDFFX1_RVT opC30_d2_reg_29_ ( .D(n3382), .SI(1'b0), .SE(n1423), .CLK(clk), 
        .QN(n1389) );
  SDFFX1_RVT opC30_d2_reg_28_ ( .D(n3382), .SI(1'b0), .SE(n1422), .CLK(clk), 
        .QN(n1387) );
  SDFFX1_RVT opC30_d2_reg_27_ ( .D(n3382), .SI(1'b0), .SE(n1421), .CLK(clk), 
        .QN(n1385) );
  SDFFX1_RVT opC30_d2_reg_26_ ( .D(n3382), .SI(1'b0), .SE(n1420), .CLK(clk), 
        .QN(n1383) );
  SDFFX1_RVT opC30_d2_reg_25_ ( .D(n3382), .SI(1'b0), .SE(n1419), .CLK(clk), 
        .QN(n1381) );
  SDFFX1_RVT opC30_d2_reg_24_ ( .D(n3382), .SI(1'b0), .SE(n1418), .CLK(clk), 
        .QN(n1379) );
  SDFFX1_RVT opC30_d2_reg_23_ ( .D(n3382), .SI(1'b0), .SE(n1417), .CLK(clk), 
        .QN(n1377) );
  SDFFX1_RVT opC30_d2_reg_22_ ( .D(n3382), .SI(1'b0), .SE(n1416), .CLK(clk), 
        .QN(n1375) );
  SDFFX1_RVT opC30_d2_reg_21_ ( .D(n3382), .SI(1'b0), .SE(n1415), .CLK(clk), 
        .QN(n1373) );
  SDFFX1_RVT opC30_d2_reg_20_ ( .D(n3382), .SI(1'b0), .SE(n1414), .CLK(clk), 
        .QN(n1371) );
  SDFFX1_RVT opC30_d2_reg_19_ ( .D(n3382), .SI(1'b0), .SE(n1413), .CLK(clk), 
        .QN(n1369) );
  SDFFX1_RVT opC30_d2_reg_18_ ( .D(n3382), .SI(1'b0), .SE(n1412), .CLK(clk), 
        .QN(n1367) );
  SDFFX1_RVT opC30_d2_reg_17_ ( .D(n3382), .SI(1'b0), .SE(n1411), .CLK(clk), 
        .QN(n1365) );
  SDFFX1_RVT opC30_d2_reg_16_ ( .D(n3381), .SI(1'b0), .SE(n1410), .CLK(clk), 
        .QN(n1363) );
  SDFFX1_RVT opC30_d2_reg_15_ ( .D(n3381), .SI(1'b0), .SE(n1409), .CLK(clk), 
        .QN(n1361) );
  SDFFX1_RVT opC30_d2_reg_14_ ( .D(n3381), .SI(1'b0), .SE(n1408), .CLK(clk), 
        .QN(n1359) );
  SDFFX1_RVT opC30_d2_reg_13_ ( .D(n3381), .SI(1'b0), .SE(n1407), .CLK(clk), 
        .QN(n1357) );
  SDFFX1_RVT opC30_d2_reg_12_ ( .D(n3381), .SI(1'b0), .SE(n1406), .CLK(clk), 
        .QN(n1355) );
  SDFFX1_RVT opC30_d2_reg_11_ ( .D(n3381), .SI(1'b0), .SE(n1405), .CLK(clk), 
        .QN(n1353) );
  SDFFX1_RVT opC30_d2_reg_10_ ( .D(n3381), .SI(1'b0), .SE(n1404), .CLK(clk), 
        .QN(n1351) );
  SDFFX1_RVT opC30_d2_reg_9_ ( .D(n3381), .SI(1'b0), .SE(n1403), .CLK(clk), 
        .QN(n1349) );
  SDFFX1_RVT opC30_d2_reg_8_ ( .D(n3381), .SI(1'b0), .SE(n1402), .CLK(clk), 
        .QN(n1347) );
  SDFFX1_RVT opC30_d2_reg_7_ ( .D(n3386), .SI(1'b0), .SE(n1401), .CLK(clk), 
        .QN(n1345) );
  SDFFX1_RVT opC30_d2_reg_6_ ( .D(n3390), .SI(1'b0), .SE(n1400), .CLK(clk), 
        .QN(n1343) );
  SDFFX1_RVT opC30_d2_reg_5_ ( .D(n3385), .SI(1'b0), .SE(n1399), .CLK(clk), 
        .QN(n1341) );
  SDFFX1_RVT opC30_d2_reg_4_ ( .D(n3381), .SI(1'b0), .SE(n1398), .CLK(clk), 
        .QN(n1339) );
  SDFFX1_RVT opC30_d2_reg_3_ ( .D(n3381), .SI(1'b0), .SE(n1397), .CLK(clk), 
        .QN(n1337) );
  SDFFX1_RVT opC30_d2_reg_2_ ( .D(n3381), .SI(1'b0), .SE(n1396), .CLK(clk), 
        .QN(n1335) );
  SDFFX1_RVT opC30_d2_reg_1_ ( .D(n3380), .SI(1'b0), .SE(n1395), .CLK(clk), 
        .QN(n1333) );
  SDFFX1_RVT opC30_d2_reg_0_ ( .D(n3380), .SI(1'b0), .SE(n1394), .CLK(clk), 
        .QN(n1331) );
  SDFFX1_RVT opC30_d1_reg_31_ ( .D(n3380), .SI(1'b0), .SE(n1393), .CLK(clk), 
        .Q(OpC30[31]) );
  SDFFX1_RVT opC30_d1_reg_30_ ( .D(n3380), .SI(1'b0), .SE(n1391), .CLK(clk), 
        .Q(OpC30[30]) );
  SDFFX1_RVT opC30_d1_reg_29_ ( .D(n3380), .SI(1'b0), .SE(n1389), .CLK(clk), 
        .Q(OpC30[29]) );
  SDFFX1_RVT opC30_d1_reg_28_ ( .D(n3380), .SI(1'b0), .SE(n1387), .CLK(clk), 
        .Q(OpC30[28]) );
  SDFFX1_RVT opC30_d1_reg_27_ ( .D(n3380), .SI(1'b0), .SE(n1385), .CLK(clk), 
        .Q(OpC30[27]) );
  SDFFX1_RVT opC30_d1_reg_26_ ( .D(n3380), .SI(1'b0), .SE(n1383), .CLK(clk), 
        .Q(OpC30[26]) );
  SDFFX1_RVT opC30_d1_reg_25_ ( .D(n3380), .SI(1'b0), .SE(n1381), .CLK(clk), 
        .Q(OpC30[25]) );
  SDFFX1_RVT opC30_d1_reg_24_ ( .D(n3380), .SI(1'b0), .SE(n1379), .CLK(clk), 
        .Q(OpC30[24]) );
  SDFFX1_RVT opC30_d1_reg_23_ ( .D(n3380), .SI(1'b0), .SE(n1377), .CLK(clk), 
        .Q(OpC30[23]) );
  SDFFX1_RVT opC30_d1_reg_22_ ( .D(n3380), .SI(1'b0), .SE(n1375), .CLK(clk), 
        .Q(OpC30[22]) );
  SDFFX1_RVT opC30_d1_reg_21_ ( .D(n3380), .SI(1'b0), .SE(n1373), .CLK(clk), 
        .Q(OpC30[21]) );
  SDFFX1_RVT opC30_d1_reg_20_ ( .D(n3380), .SI(1'b0), .SE(n1371), .CLK(clk), 
        .Q(OpC30[20]) );
  SDFFX1_RVT opC30_d1_reg_19_ ( .D(n3379), .SI(1'b0), .SE(n1369), .CLK(clk), 
        .Q(OpC30[19]) );
  SDFFX1_RVT opC30_d1_reg_18_ ( .D(n3379), .SI(1'b0), .SE(n1367), .CLK(clk), 
        .Q(OpC30[18]) );
  SDFFX1_RVT opC30_d1_reg_17_ ( .D(n3379), .SI(1'b0), .SE(n1365), .CLK(clk), 
        .Q(OpC30[17]) );
  SDFFX1_RVT opC30_d1_reg_16_ ( .D(n3379), .SI(1'b0), .SE(n1363), .CLK(clk), 
        .Q(OpC30[16]) );
  SDFFX1_RVT opC30_d1_reg_15_ ( .D(n3379), .SI(1'b0), .SE(n1361), .CLK(clk), 
        .Q(OpC30[15]) );
  SDFFX1_RVT opC30_d1_reg_14_ ( .D(n3379), .SI(1'b0), .SE(n1359), .CLK(clk), 
        .Q(OpC30[14]) );
  SDFFX1_RVT opC30_d1_reg_13_ ( .D(n3379), .SI(1'b0), .SE(n1357), .CLK(clk), 
        .Q(OpC30[13]) );
  SDFFX1_RVT opC30_d1_reg_12_ ( .D(n3379), .SI(1'b0), .SE(n1355), .CLK(clk), 
        .Q(OpC30[12]) );
  SDFFX1_RVT opC30_d1_reg_11_ ( .D(n3379), .SI(1'b0), .SE(n1353), .CLK(clk), 
        .Q(OpC30[11]) );
  SDFFX1_RVT opC30_d1_reg_10_ ( .D(n3379), .SI(1'b0), .SE(n1351), .CLK(clk), 
        .Q(OpC30[10]) );
  SDFFX1_RVT opC30_d1_reg_9_ ( .D(n3379), .SI(1'b0), .SE(n1349), .CLK(clk), 
        .Q(OpC30[9]) );
  SDFFX1_RVT opC30_d1_reg_8_ ( .D(n3379), .SI(1'b0), .SE(n1347), .CLK(clk), 
        .Q(OpC30[8]) );
  SDFFX1_RVT opC30_d1_reg_7_ ( .D(n3379), .SI(1'b0), .SE(n1345), .CLK(clk), 
        .Q(OpC30[7]) );
  SDFFX1_RVT opC30_d1_reg_6_ ( .D(n3379), .SI(1'b0), .SE(n1343), .CLK(clk), 
        .Q(OpC30[6]) );
  SDFFX1_RVT opC30_d1_reg_5_ ( .D(n3378), .SI(1'b0), .SE(n1341), .CLK(clk), 
        .Q(OpC30[5]) );
  SDFFX1_RVT opC30_d1_reg_4_ ( .D(n3378), .SI(1'b0), .SE(n1339), .CLK(clk), 
        .Q(OpC30[4]) );
  SDFFX1_RVT opC30_d1_reg_3_ ( .D(n3378), .SI(1'b0), .SE(n1337), .CLK(clk), 
        .Q(OpC30[3]) );
  SDFFX1_RVT opC30_d1_reg_2_ ( .D(n3378), .SI(1'b0), .SE(n1335), .CLK(clk), 
        .Q(OpC30[2]) );
  SDFFX1_RVT opC30_d1_reg_1_ ( .D(n3378), .SI(1'b0), .SE(n1333), .CLK(clk), 
        .Q(OpC30[1]) );
  SDFFX1_RVT opC30_d1_reg_0_ ( .D(n3378), .SI(1'b0), .SE(n1331), .CLK(clk), 
        .Q(OpC30[0]) );
  SDFFX1_RVT opC13_d1_reg_31_ ( .D(n3378), .SI(1'b0), .SE(n1297), .CLK(clk), 
        .Q(OpC13[31]) );
  SDFFX1_RVT opC13_d1_reg_30_ ( .D(n3378), .SI(1'b0), .SE(n1296), .CLK(clk), 
        .Q(OpC13[30]) );
  SDFFX1_RVT opC13_d1_reg_29_ ( .D(n3378), .SI(1'b0), .SE(n1295), .CLK(clk), 
        .Q(OpC13[29]) );
  SDFFX1_RVT opC13_d1_reg_28_ ( .D(n3378), .SI(1'b0), .SE(n1294), .CLK(clk), 
        .Q(OpC13[28]) );
  SDFFX1_RVT opC13_d1_reg_27_ ( .D(n3378), .SI(1'b0), .SE(n1293), .CLK(clk), 
        .Q(OpC13[27]) );
  SDFFX1_RVT opC13_d1_reg_26_ ( .D(n3378), .SI(1'b0), .SE(n1292), .CLK(clk), 
        .Q(OpC13[26]) );
  SDFFX1_RVT opC13_d1_reg_25_ ( .D(n3378), .SI(1'b0), .SE(n1291), .CLK(clk), 
        .Q(OpC13[25]) );
  SDFFX1_RVT opC13_d1_reg_24_ ( .D(n3378), .SI(1'b0), .SE(n1290), .CLK(clk), 
        .Q(OpC13[24]) );
  SDFFX1_RVT opC13_d1_reg_23_ ( .D(n3377), .SI(1'b0), .SE(n1289), .CLK(clk), 
        .Q(OpC13[23]) );
  SDFFX1_RVT opC13_d1_reg_22_ ( .D(n3377), .SI(1'b0), .SE(n1288), .CLK(clk), 
        .Q(OpC13[22]) );
  SDFFX1_RVT opC13_d1_reg_21_ ( .D(n3377), .SI(1'b0), .SE(n1287), .CLK(clk), 
        .Q(OpC13[21]) );
  SDFFX1_RVT opC13_d1_reg_20_ ( .D(n3377), .SI(1'b0), .SE(n1286), .CLK(clk), 
        .Q(OpC13[20]) );
  SDFFX1_RVT opC13_d1_reg_19_ ( .D(n3377), .SI(1'b0), .SE(n1285), .CLK(clk), 
        .Q(OpC13[19]) );
  SDFFX1_RVT opC13_d1_reg_18_ ( .D(n3377), .SI(1'b0), .SE(n1284), .CLK(clk), 
        .Q(OpC13[18]) );
  SDFFX1_RVT opC13_d1_reg_17_ ( .D(n3377), .SI(1'b0), .SE(n1283), .CLK(clk), 
        .Q(OpC13[17]) );
  SDFFX1_RVT opC13_d1_reg_16_ ( .D(n3377), .SI(1'b0), .SE(n1282), .CLK(clk), 
        .Q(OpC13[16]) );
  SDFFX1_RVT opC13_d1_reg_15_ ( .D(n3377), .SI(1'b0), .SE(n1281), .CLK(clk), 
        .Q(OpC13[15]) );
  SDFFX1_RVT opC13_d1_reg_14_ ( .D(n3377), .SI(1'b0), .SE(n1280), .CLK(clk), 
        .Q(OpC13[14]) );
  SDFFX1_RVT opC13_d1_reg_13_ ( .D(n3377), .SI(1'b0), .SE(n1279), .CLK(clk), 
        .Q(OpC13[13]) );
  SDFFX1_RVT opC13_d1_reg_12_ ( .D(n3377), .SI(1'b0), .SE(n1278), .CLK(clk), 
        .Q(OpC13[12]) );
  SDFFX1_RVT opC13_d1_reg_11_ ( .D(n3377), .SI(1'b0), .SE(n1277), .CLK(clk), 
        .Q(OpC13[11]) );
  SDFFX1_RVT opC13_d1_reg_10_ ( .D(n3377), .SI(1'b0), .SE(n1276), .CLK(clk), 
        .Q(OpC13[10]) );
  SDFFX1_RVT opC13_d1_reg_9_ ( .D(n3376), .SI(1'b0), .SE(n1275), .CLK(clk), 
        .Q(OpC13[9]) );
  SDFFX1_RVT opC13_d1_reg_8_ ( .D(n3376), .SI(1'b0), .SE(n1274), .CLK(clk), 
        .Q(OpC13[8]) );
  SDFFX1_RVT opC13_d1_reg_7_ ( .D(n3376), .SI(1'b0), .SE(n1273), .CLK(clk), 
        .Q(OpC13[7]) );
  SDFFX1_RVT opC13_d1_reg_6_ ( .D(n3376), .SI(1'b0), .SE(n1272), .CLK(clk), 
        .Q(OpC13[6]) );
  SDFFX1_RVT opC13_d1_reg_5_ ( .D(n3376), .SI(1'b0), .SE(n1271), .CLK(clk), 
        .Q(OpC13[5]) );
  SDFFX1_RVT opC13_d1_reg_4_ ( .D(n3376), .SI(1'b0), .SE(n1270), .CLK(clk), 
        .Q(OpC13[4]) );
  SDFFX1_RVT opC13_d1_reg_3_ ( .D(n3376), .SI(1'b0), .SE(n1269), .CLK(clk), 
        .Q(OpC13[3]) );
  SDFFX1_RVT opC13_d1_reg_2_ ( .D(n3376), .SI(1'b0), .SE(n1268), .CLK(clk), 
        .Q(OpC13[2]) );
  SDFFX1_RVT opC13_d1_reg_1_ ( .D(n3376), .SI(1'b0), .SE(n1267), .CLK(clk), 
        .Q(OpC13[1]) );
  SDFFX1_RVT opC13_d1_reg_0_ ( .D(n3376), .SI(1'b0), .SE(n1266), .CLK(clk), 
        .Q(OpC13[0]) );
  SDFFX1_RVT opC22_d1_reg_31_ ( .D(n3376), .SI(1'b0), .SE(n1233), .CLK(clk), 
        .Q(OpC22[31]) );
  SDFFX1_RVT opC22_d1_reg_30_ ( .D(n3376), .SI(1'b0), .SE(n1232), .CLK(clk), 
        .Q(OpC22[30]) );
  SDFFX1_RVT opC22_d1_reg_29_ ( .D(n3375), .SI(1'b0), .SE(n1231), .CLK(clk), 
        .Q(OpC22[29]) );
  SDFFX1_RVT opC22_d1_reg_28_ ( .D(n3375), .SI(1'b0), .SE(n1230), .CLK(clk), 
        .Q(OpC22[28]) );
  SDFFX1_RVT opC22_d1_reg_27_ ( .D(n3375), .SI(1'b0), .SE(n1229), .CLK(clk), 
        .Q(OpC22[27]) );
  SDFFX1_RVT opC22_d1_reg_26_ ( .D(n3375), .SI(1'b0), .SE(n1228), .CLK(clk), 
        .Q(OpC22[26]) );
  SDFFX1_RVT opC22_d1_reg_25_ ( .D(n3375), .SI(1'b0), .SE(n1227), .CLK(clk), 
        .Q(OpC22[25]) );
  SDFFX1_RVT opC22_d1_reg_24_ ( .D(n3375), .SI(1'b0), .SE(n1226), .CLK(clk), 
        .Q(OpC22[24]) );
  SDFFX1_RVT opC22_d1_reg_23_ ( .D(n3375), .SI(1'b0), .SE(n1225), .CLK(clk), 
        .Q(OpC22[23]) );
  SDFFX1_RVT opC22_d1_reg_22_ ( .D(n3375), .SI(1'b0), .SE(n1224), .CLK(clk), 
        .Q(OpC22[22]) );
  SDFFX1_RVT opC22_d1_reg_21_ ( .D(n3375), .SI(1'b0), .SE(n1223), .CLK(clk), 
        .Q(OpC22[21]) );
  SDFFX1_RVT opC22_d1_reg_20_ ( .D(n3375), .SI(1'b0), .SE(n1222), .CLK(clk), 
        .Q(OpC22[20]) );
  SDFFX1_RVT opC22_d1_reg_19_ ( .D(n3375), .SI(1'b0), .SE(n1221), .CLK(clk), 
        .Q(OpC22[19]) );
  SDFFX1_RVT opC22_d1_reg_18_ ( .D(n3375), .SI(1'b0), .SE(n1220), .CLK(clk), 
        .Q(OpC22[18]) );
  SDFFX1_RVT opC22_d1_reg_17_ ( .D(n3375), .SI(1'b0), .SE(n1219), .CLK(clk), 
        .Q(OpC22[17]) );
  SDFFX1_RVT opC22_d1_reg_16_ ( .D(n3375), .SI(1'b0), .SE(n1218), .CLK(clk), 
        .Q(OpC22[16]) );
  SDFFX1_RVT opC22_d1_reg_15_ ( .D(n3374), .SI(1'b0), .SE(n1217), .CLK(clk), 
        .Q(OpC22[15]) );
  SDFFX1_RVT opC22_d1_reg_14_ ( .D(n3374), .SI(1'b0), .SE(n1216), .CLK(clk), 
        .Q(OpC22[14]) );
  SDFFX1_RVT opC22_d1_reg_13_ ( .D(n3374), .SI(1'b0), .SE(n1215), .CLK(clk), 
        .Q(OpC22[13]) );
  SDFFX1_RVT opC22_d1_reg_12_ ( .D(n3374), .SI(1'b0), .SE(n1214), .CLK(clk), 
        .Q(OpC22[12]) );
  SDFFX1_RVT opC22_d1_reg_11_ ( .D(n3374), .SI(1'b0), .SE(n1213), .CLK(clk), 
        .Q(OpC22[11]) );
  SDFFX1_RVT opC22_d1_reg_10_ ( .D(n3374), .SI(1'b0), .SE(n1212), .CLK(clk), 
        .Q(OpC22[10]) );
  SDFFX1_RVT opC22_d1_reg_9_ ( .D(n3374), .SI(1'b0), .SE(n1211), .CLK(clk), 
        .Q(OpC22[9]) );
  SDFFX1_RVT opC22_d1_reg_8_ ( .D(n3374), .SI(1'b0), .SE(n1210), .CLK(clk), 
        .Q(OpC22[8]) );
  SDFFX1_RVT opC22_d1_reg_7_ ( .D(n3376), .SI(1'b0), .SE(n1209), .CLK(clk), 
        .Q(OpC22[7]) );
  SDFFX1_RVT opC22_d1_reg_6_ ( .D(n3374), .SI(1'b0), .SE(n1208), .CLK(clk), 
        .Q(OpC22[6]) );
  SDFFX1_RVT opC22_d1_reg_5_ ( .D(n3374), .SI(1'b0), .SE(n1207), .CLK(clk), 
        .Q(OpC22[5]) );
  SDFFX1_RVT opC22_d1_reg_4_ ( .D(n3374), .SI(1'b0), .SE(n1206), .CLK(clk), 
        .Q(OpC22[4]) );
  SDFFX1_RVT opC22_d1_reg_3_ ( .D(n3374), .SI(1'b0), .SE(n1205), .CLK(clk), 
        .Q(OpC22[3]) );
  SDFFX1_RVT opC22_d1_reg_2_ ( .D(n3374), .SI(1'b0), .SE(n1204), .CLK(clk), 
        .Q(OpC22[2]) );
  SDFFX1_RVT opC22_d1_reg_1_ ( .D(n3374), .SI(1'b0), .SE(n1203), .CLK(clk), 
        .Q(OpC22[1]) );
  SDFFX1_RVT opC22_d1_reg_0_ ( .D(n3373), .SI(1'b0), .SE(n1202), .CLK(clk), 
        .Q(OpC22[0]) );
  SDFFX1_RVT opC31_d1_reg_31_ ( .D(n3373), .SI(1'b0), .SE(n1169), .CLK(clk), 
        .Q(OpC31[31]) );
  SDFFX1_RVT opC31_d1_reg_30_ ( .D(n3373), .SI(1'b0), .SE(n1167), .CLK(clk), 
        .Q(OpC31[30]) );
  SDFFX1_RVT opC31_d1_reg_29_ ( .D(n3373), .SI(1'b0), .SE(n1165), .CLK(clk), 
        .Q(OpC31[29]) );
  SDFFX1_RVT opC31_d1_reg_28_ ( .D(n3373), .SI(1'b0), .SE(n1163), .CLK(clk), 
        .Q(OpC31[28]) );
  SDFFX1_RVT opC31_d1_reg_27_ ( .D(n3373), .SI(1'b0), .SE(n1161), .CLK(clk), 
        .Q(OpC31[27]) );
  SDFFX1_RVT opC31_d1_reg_26_ ( .D(n3373), .SI(1'b0), .SE(n1159), .CLK(clk), 
        .Q(OpC31[26]) );
  SDFFX1_RVT opC31_d1_reg_25_ ( .D(n3373), .SI(1'b0), .SE(n1157), .CLK(clk), 
        .Q(OpC31[25]) );
  SDFFX1_RVT opC31_d1_reg_24_ ( .D(n3373), .SI(1'b0), .SE(n1155), .CLK(clk), 
        .Q(OpC31[24]) );
  SDFFX1_RVT opC31_d1_reg_23_ ( .D(n3373), .SI(1'b0), .SE(n1153), .CLK(clk), 
        .Q(OpC31[23]) );
  SDFFX1_RVT opC31_d1_reg_22_ ( .D(n3373), .SI(1'b0), .SE(n1151), .CLK(clk), 
        .Q(OpC31[22]) );
  SDFFX1_RVT opC31_d1_reg_21_ ( .D(n3373), .SI(1'b0), .SE(n1149), .CLK(clk), 
        .Q(OpC31[21]) );
  SDFFX1_RVT opC31_d1_reg_20_ ( .D(n3373), .SI(1'b0), .SE(n1147), .CLK(clk), 
        .Q(OpC31[20]) );
  SDFFX1_RVT opC31_d1_reg_19_ ( .D(n3373), .SI(1'b0), .SE(n1145), .CLK(clk), 
        .Q(OpC31[19]) );
  SDFFX1_RVT opC31_d1_reg_18_ ( .D(n3466), .SI(1'b0), .SE(n1143), .CLK(clk), 
        .Q(OpC31[18]) );
  SDFFX1_RVT opC31_d1_reg_17_ ( .D(n3466), .SI(1'b0), .SE(n1141), .CLK(clk), 
        .Q(OpC31[17]) );
  SDFFX1_RVT opC31_d1_reg_16_ ( .D(n3466), .SI(1'b0), .SE(n1139), .CLK(clk), 
        .Q(OpC31[16]) );
  SDFFX1_RVT opC31_d1_reg_15_ ( .D(n3466), .SI(1'b0), .SE(n1137), .CLK(clk), 
        .Q(OpC31[15]) );
  SDFFX1_RVT opC31_d1_reg_14_ ( .D(n3408), .SI(1'b0), .SE(n1135), .CLK(clk), 
        .Q(OpC31[14]) );
  SDFFX1_RVT opC31_d1_reg_13_ ( .D(n3465), .SI(1'b0), .SE(n1133), .CLK(clk), 
        .Q(OpC31[13]) );
  SDFFX1_RVT opC31_d1_reg_12_ ( .D(n3346), .SI(1'b0), .SE(n1131), .CLK(clk), 
        .Q(OpC31[12]) );
  SDFFX1_RVT opC31_d1_reg_11_ ( .D(n3477), .SI(1'b0), .SE(n1129), .CLK(clk), 
        .Q(OpC31[11]) );
  SDFFX1_RVT opC31_d1_reg_10_ ( .D(n3479), .SI(1'b0), .SE(n1127), .CLK(clk), 
        .Q(OpC31[10]) );
  SDFFX1_RVT opC31_d1_reg_9_ ( .D(n3478), .SI(1'b0), .SE(n1125), .CLK(clk), 
        .Q(OpC31[9]) );
  SDFFX1_RVT opC31_d1_reg_8_ ( .D(n3480), .SI(1'b0), .SE(n1123), .CLK(clk), 
        .Q(OpC31[8]) );
  SDFFX1_RVT opC31_d1_reg_7_ ( .D(n3444), .SI(1'b0), .SE(n1121), .CLK(clk), 
        .Q(OpC31[7]) );
  SDFFX1_RVT opC31_d1_reg_6_ ( .D(n3443), .SI(1'b0), .SE(n1119), .CLK(clk), 
        .Q(OpC31[6]) );
  SDFFX1_RVT opC31_d1_reg_5_ ( .D(n3464), .SI(1'b0), .SE(n1117), .CLK(clk), 
        .Q(OpC31[5]) );
  SDFFX1_RVT opC31_d1_reg_4_ ( .D(n3481), .SI(1'b0), .SE(n1115), .CLK(clk), 
        .Q(OpC31[4]) );
  SDFFX1_RVT opC31_d1_reg_2_ ( .D(n3376), .SI(1'b0), .SE(n1111), .CLK(clk), 
        .Q(OpC31[2]) );
  SDFFX1_RVT opC31_d1_reg_1_ ( .D(n3381), .SI(1'b0), .SE(n1109), .CLK(clk), 
        .Q(OpC31[1]) );
  SDFFX1_RVT opC31_d1_reg_0_ ( .D(n3413), .SI(1'b0), .SE(n1107), .CLK(clk), 
        .Q(OpC31[0]) );
  AO22X1_RVT U3 ( .A1(n3573), .A2(BankAddr[9]), .A3(N25), .A4(n2), .Y(n3216)
         );
  AO22X1_RVT U4 ( .A1(n3573), .A2(BankAddr[8]), .A3(N24), .A4(n2), .Y(n3217)
         );
  AO22X1_RVT U5 ( .A1(n3573), .A2(BankAddr[7]), .A3(N23), .A4(n2), .Y(n3218)
         );
  AO22X1_RVT U6 ( .A1(n3573), .A2(BankAddr[6]), .A3(N22), .A4(n2), .Y(n3219)
         );
  AO22X1_RVT U7 ( .A1(n3573), .A2(BankAddr[5]), .A3(N21), .A4(n2), .Y(n3220)
         );
  AO22X1_RVT U8 ( .A1(n3573), .A2(BankAddr[4]), .A3(N20), .A4(n2), .Y(n3221)
         );
  AO22X1_RVT U9 ( .A1(n3573), .A2(BankAddr[3]), .A3(N19), .A4(n2), .Y(n3222)
         );
  AO22X1_RVT U10 ( .A1(n3573), .A2(BankAddr[2]), .A3(N18), .A4(n2), .Y(n3223)
         );
  AO22X1_RVT U11 ( .A1(n3573), .A2(BankAddr[1]), .A3(N17), .A4(n2), .Y(n3224)
         );
  AO22X1_RVT U12 ( .A1(n3573), .A2(BankAddr[0]), .A3(N16), .A4(n2), .Y(n3225)
         );
  AND2X1_RVT U13 ( .A1(rstnAddr), .A2(n3), .Y(n2) );
  NAND2X0_RVT U15 ( .A1(n3574), .A2(rstnAddr), .Y(n3) );
  AO22X1_RVT U17 ( .A1(n3441), .A2(opC00_out[0]), .A3(n1042), .A4(n3569), .Y(
        n3184) );
  AO22X1_RVT U18 ( .A1(opC00_out[1]), .A2(n3468), .A3(n1043), .A4(n3569), .Y(
        n3185) );
  AO22X1_RVT U19 ( .A1(opC00_out[2]), .A2(n3372), .A3(n1044), .A4(n3569), .Y(
        n3186) );
  AO22X1_RVT U20 ( .A1(opC00_out[3]), .A2(n3372), .A3(n1045), .A4(n3569), .Y(
        n3187) );
  AO22X1_RVT U21 ( .A1(opC00_out[4]), .A2(n3457), .A3(n1046), .A4(n3569), .Y(
        n3188) );
  AO22X1_RVT U22 ( .A1(opC00_out[5]), .A2(n3463), .A3(n1047), .A4(n3569), .Y(
        n3189) );
  AO22X1_RVT U23 ( .A1(opC00_out[6]), .A2(n3461), .A3(n1048), .A4(n3569), .Y(
        n3190) );
  AO22X1_RVT U24 ( .A1(opC00_out[7]), .A2(n3462), .A3(n1049), .A4(n3568), .Y(
        n3191) );
  AO22X1_RVT U25 ( .A1(opC00_out[8]), .A2(n3474), .A3(n1050), .A4(n3568), .Y(
        n3192) );
  AO22X1_RVT U26 ( .A1(opC00_out[9]), .A2(n3464), .A3(n1051), .A4(n3568), .Y(
        n3193) );
  AO22X1_RVT U27 ( .A1(opC00_out[10]), .A2(n3455), .A3(n1052), .A4(n3568), .Y(
        n3194) );
  AO22X1_RVT U28 ( .A1(opC00_out[11]), .A2(n3457), .A3(n1053), .A4(n3568), .Y(
        n3195) );
  AO22X1_RVT U29 ( .A1(opC00_out[12]), .A2(n3475), .A3(n1054), .A4(n3568), .Y(
        n3196) );
  AO22X1_RVT U30 ( .A1(opC00_out[13]), .A2(n3476), .A3(n1055), .A4(n3568), .Y(
        n3197) );
  AO22X1_RVT U31 ( .A1(opC00_out[14]), .A2(n3372), .A3(n1056), .A4(n3568), .Y(
        n3198) );
  AO22X1_RVT U32 ( .A1(opC00_out[15]), .A2(n3372), .A3(n1057), .A4(n3568), .Y(
        n3199) );
  AO22X1_RVT U33 ( .A1(opC00_out[16]), .A2(n3455), .A3(n1058), .A4(n3568), .Y(
        n3200) );
  AO22X1_RVT U34 ( .A1(opC00_out[17]), .A2(n3372), .A3(n1059), .A4(n3568), .Y(
        n3201) );
  AO22X1_RVT U35 ( .A1(opC00_out[18]), .A2(n3372), .A3(n1060), .A4(n3568), .Y(
        n3202) );
  AO22X1_RVT U36 ( .A1(opC00_out[19]), .A2(n3372), .A3(n1061), .A4(n3568), .Y(
        n3203) );
  AO22X1_RVT U37 ( .A1(opC00_out[20]), .A2(n3372), .A3(n1062), .A4(n3567), .Y(
        n3204) );
  AO22X1_RVT U38 ( .A1(opC00_out[21]), .A2(n3372), .A3(n1063), .A4(n3567), .Y(
        n3205) );
  AO22X1_RVT U39 ( .A1(opC00_out[22]), .A2(n3372), .A3(n1064), .A4(n3567), .Y(
        n3206) );
  AO22X1_RVT U40 ( .A1(opC00_out[23]), .A2(n3372), .A3(n1065), .A4(n3567), .Y(
        n3207) );
  AO22X1_RVT U41 ( .A1(opC00_out[24]), .A2(n3372), .A3(n1066), .A4(n3567), .Y(
        n3208) );
  AO22X1_RVT U42 ( .A1(opC00_out[25]), .A2(n3464), .A3(n1067), .A4(n3567), .Y(
        n3209) );
  AO22X1_RVT U43 ( .A1(opC00_out[26]), .A2(n3372), .A3(n1068), .A4(n3567), .Y(
        n3210) );
  AO22X1_RVT U44 ( .A1(opC00_out[27]), .A2(n3464), .A3(n1069), .A4(n3567), .Y(
        n3211) );
  AO22X1_RVT U45 ( .A1(opC00_out[28]), .A2(n3464), .A3(n1070), .A4(n3567), .Y(
        n3212) );
  AO22X1_RVT U46 ( .A1(opC00_out[29]), .A2(n3464), .A3(n1071), .A4(n3567), .Y(
        n3213) );
  AO22X1_RVT U47 ( .A1(opC00_out[30]), .A2(n3367), .A3(n1072), .A4(n3567), .Y(
        n3214) );
  AO22X1_RVT U48 ( .A1(opC00_out[31]), .A2(n3367), .A3(n1073), .A4(n3567), .Y(
        n3215) );
  OR3X1_RVT U50 ( .A1(n6), .A2(n7), .A3(n8), .Y(ipB3[9]) );
  AO221X1_RVT U51 ( .A1(MemOutputB3[9]), .A2(n3299), .A3(MemOutputB3[41]), 
        .A4(n3545), .A5(n11), .Y(n8) );
  AO22X1_RVT U52 ( .A1(MemOutputB3[73]), .A2(n3525), .A3(MemOutputB3[105]), 
        .A4(n3506), .Y(n11) );
  AO22X1_RVT U53 ( .A1(MemOutputB3[169]), .A2(n3264), .A3(MemOutputB3[137]), 
        .A4(n3273), .Y(n7) );
  AO22X1_RVT U54 ( .A1(MemOutputB3[201]), .A2(n3484), .A3(MemOutputB3[233]), 
        .A4(n3334), .Y(n6) );
  OR3X1_RVT U55 ( .A1(n18), .A2(n19), .A3(n20), .Y(ipB3[8]) );
  AO221X1_RVT U56 ( .A1(MemOutputB3[8]), .A2(n3298), .A3(MemOutputB3[40]), 
        .A4(n3545), .A5(n21), .Y(n20) );
  AO22X1_RVT U57 ( .A1(MemOutputB3[72]), .A2(n3525), .A3(MemOutputB3[104]), 
        .A4(n3506), .Y(n21) );
  AO22X1_RVT U58 ( .A1(MemOutputB3[168]), .A2(n3265), .A3(MemOutputB3[136]), 
        .A4(n3281), .Y(n19) );
  AO22X1_RVT U59 ( .A1(MemOutputB3[200]), .A2(n3484), .A3(MemOutputB3[232]), 
        .A4(n3333), .Y(n18) );
  OR3X1_RVT U60 ( .A1(n22), .A2(n23), .A3(n24), .Y(ipB3[7]) );
  AO221X1_RVT U61 ( .A1(MemOutputB3[7]), .A2(n3298), .A3(MemOutputB3[39]), 
        .A4(n3545), .A5(n25), .Y(n24) );
  AO22X1_RVT U62 ( .A1(MemOutputB3[71]), .A2(n3525), .A3(MemOutputB3[103]), 
        .A4(n3506), .Y(n25) );
  AO22X1_RVT U63 ( .A1(MemOutputB3[167]), .A2(n3249), .A3(MemOutputB3[135]), 
        .A4(n3276), .Y(n23) );
  AO22X1_RVT U64 ( .A1(MemOutputB3[199]), .A2(n3484), .A3(MemOutputB3[231]), 
        .A4(n3324), .Y(n22) );
  OR3X1_RVT U65 ( .A1(n26), .A2(n27), .A3(n28), .Y(ipB3[6]) );
  AO221X1_RVT U66 ( .A1(MemOutputB3[6]), .A2(n3297), .A3(MemOutputB3[38]), 
        .A4(n3545), .A5(n29), .Y(n28) );
  AO22X1_RVT U67 ( .A1(MemOutputB3[70]), .A2(n3525), .A3(MemOutputB3[102]), 
        .A4(n3506), .Y(n29) );
  AO22X1_RVT U68 ( .A1(MemOutputB3[166]), .A2(n3249), .A3(MemOutputB3[134]), 
        .A4(n454), .Y(n27) );
  AO22X1_RVT U69 ( .A1(MemOutputB3[198]), .A2(n3484), .A3(MemOutputB3[230]), 
        .A4(n3336), .Y(n26) );
  OR3X1_RVT U70 ( .A1(n30), .A2(n31), .A3(n32), .Y(ipB3[5]) );
  AO221X1_RVT U71 ( .A1(MemOutputB3[5]), .A2(n3297), .A3(MemOutputB3[37]), 
        .A4(n3545), .A5(n33), .Y(n32) );
  AO22X1_RVT U72 ( .A1(MemOutputB3[69]), .A2(n3525), .A3(MemOutputB3[101]), 
        .A4(n3506), .Y(n33) );
  AO22X1_RVT U73 ( .A1(MemOutputB3[165]), .A2(n3247), .A3(MemOutputB3[133]), 
        .A4(n506), .Y(n31) );
  AO22X1_RVT U74 ( .A1(MemOutputB3[197]), .A2(n3484), .A3(MemOutputB3[229]), 
        .A4(n3326), .Y(n30) );
  OR3X1_RVT U75 ( .A1(n34), .A2(n35), .A3(n36), .Y(ipB3[4]) );
  AO221X1_RVT U76 ( .A1(MemOutputB3[4]), .A2(n3296), .A3(MemOutputB3[36]), 
        .A4(n3545), .A5(n37), .Y(n36) );
  AO22X1_RVT U77 ( .A1(MemOutputB3[68]), .A2(n3525), .A3(MemOutputB3[100]), 
        .A4(n3506), .Y(n37) );
  AO22X1_RVT U78 ( .A1(MemOutputB3[164]), .A2(n3247), .A3(MemOutputB3[132]), 
        .A4(n506), .Y(n35) );
  AO22X1_RVT U79 ( .A1(MemOutputB3[196]), .A2(n3484), .A3(MemOutputB3[228]), 
        .A4(n3336), .Y(n34) );
  OR3X1_RVT U80 ( .A1(n38), .A2(n39), .A3(n40), .Y(ipB3[3]) );
  AO221X1_RVT U81 ( .A1(MemOutputB3[3]), .A2(n3297), .A3(MemOutputB3[35]), 
        .A4(n3545), .A5(n41), .Y(n40) );
  AO22X1_RVT U82 ( .A1(MemOutputB3[67]), .A2(n3525), .A3(MemOutputB3[99]), 
        .A4(n3506), .Y(n41) );
  AO22X1_RVT U83 ( .A1(MemOutputB3[163]), .A2(n3248), .A3(MemOutputB3[131]), 
        .A4(n3270), .Y(n39) );
  AO22X1_RVT U84 ( .A1(MemOutputB3[195]), .A2(n3484), .A3(MemOutputB3[227]), 
        .A4(n3326), .Y(n38) );
  OR3X1_RVT U85 ( .A1(n42), .A2(n43), .A3(n44), .Y(ipB3[31]) );
  AO221X1_RVT U86 ( .A1(MemOutputB3[31]), .A2(n3296), .A3(MemOutputB3[63]), 
        .A4(n3545), .A5(n45), .Y(n44) );
  AO22X1_RVT U87 ( .A1(MemOutputB3[95]), .A2(n3525), .A3(MemOutputB3[127]), 
        .A4(n3506), .Y(n45) );
  AO22X1_RVT U88 ( .A1(MemOutputB3[191]), .A2(n3264), .A3(MemOutputB3[159]), 
        .A4(n3283), .Y(n43) );
  AO22X1_RVT U89 ( .A1(MemOutputB3[223]), .A2(n3484), .A3(MemOutputB3[255]), 
        .A4(n3325), .Y(n42) );
  OR3X1_RVT U90 ( .A1(n46), .A2(n47), .A3(n48), .Y(ipB3[30]) );
  AO221X1_RVT U91 ( .A1(MemOutputB3[30]), .A2(n3298), .A3(MemOutputB3[62]), 
        .A4(n3545), .A5(n49), .Y(n48) );
  AO22X1_RVT U92 ( .A1(MemOutputB3[94]), .A2(n3525), .A3(MemOutputB3[126]), 
        .A4(n3506), .Y(n49) );
  AO22X1_RVT U93 ( .A1(MemOutputB3[190]), .A2(n514), .A3(MemOutputB3[158]), 
        .A4(n3272), .Y(n47) );
  AO22X1_RVT U94 ( .A1(MemOutputB3[222]), .A2(n3484), .A3(MemOutputB3[254]), 
        .A4(n3333), .Y(n46) );
  OR3X1_RVT U95 ( .A1(n50), .A2(n51), .A3(n52), .Y(ipB3[2]) );
  AO221X1_RVT U96 ( .A1(MemOutputB3[2]), .A2(n3298), .A3(MemOutputB3[34]), 
        .A4(n3545), .A5(n53), .Y(n52) );
  AO22X1_RVT U97 ( .A1(MemOutputB3[66]), .A2(n3525), .A3(MemOutputB3[98]), 
        .A4(n3506), .Y(n53) );
  AO22X1_RVT U98 ( .A1(MemOutputB3[162]), .A2(n3263), .A3(MemOutputB3[130]), 
        .A4(n3277), .Y(n51) );
  AO22X1_RVT U99 ( .A1(MemOutputB3[194]), .A2(n3484), .A3(MemOutputB3[226]), 
        .A4(n3323), .Y(n50) );
  OR3X1_RVT U100 ( .A1(n54), .A2(n55), .A3(n56), .Y(ipB3[29]) );
  AO221X1_RVT U101 ( .A1(MemOutputB3[29]), .A2(n3296), .A3(MemOutputB3[61]), 
        .A4(n3545), .A5(n57), .Y(n56) );
  AO22X1_RVT U102 ( .A1(MemOutputB3[93]), .A2(n3525), .A3(MemOutputB3[125]), 
        .A4(n3506), .Y(n57) );
  AO22X1_RVT U103 ( .A1(MemOutputB3[189]), .A2(n3264), .A3(MemOutputB3[157]), 
        .A4(n452), .Y(n55) );
  AO22X1_RVT U104 ( .A1(MemOutputB3[221]), .A2(n3484), .A3(MemOutputB3[253]), 
        .A4(n3323), .Y(n54) );
  OR3X1_RVT U105 ( .A1(n58), .A2(n59), .A3(n60), .Y(ipB3[28]) );
  AO221X1_RVT U106 ( .A1(MemOutputB3[28]), .A2(n3304), .A3(MemOutputB3[60]), 
        .A4(n3545), .A5(n61), .Y(n60) );
  AO22X1_RVT U107 ( .A1(MemOutputB3[92]), .A2(n3525), .A3(MemOutputB3[124]), 
        .A4(n3506), .Y(n61) );
  AO22X1_RVT U108 ( .A1(MemOutputB3[188]), .A2(n3263), .A3(MemOutputB3[156]), 
        .A4(n3282), .Y(n59) );
  AO22X1_RVT U109 ( .A1(MemOutputB3[220]), .A2(n3484), .A3(MemOutputB3[252]), 
        .A4(n3336), .Y(n58) );
  OR3X1_RVT U110 ( .A1(n62), .A2(n63), .A3(n64), .Y(ipB3[27]) );
  AO221X1_RVT U111 ( .A1(MemOutputB3[27]), .A2(n3298), .A3(MemOutputB3[59]), 
        .A4(n3546), .A5(n65), .Y(n64) );
  AO22X1_RVT U112 ( .A1(MemOutputB3[91]), .A2(n3526), .A3(MemOutputB3[123]), 
        .A4(n3507), .Y(n65) );
  AO22X1_RVT U113 ( .A1(MemOutputB3[187]), .A2(n3265), .A3(MemOutputB3[155]), 
        .A4(n3283), .Y(n63) );
  AO22X1_RVT U114 ( .A1(MemOutputB3[219]), .A2(n3485), .A3(MemOutputB3[251]), 
        .A4(n3323), .Y(n62) );
  OR3X1_RVT U115 ( .A1(n66), .A2(n67), .A3(n68), .Y(ipB3[26]) );
  AO221X1_RVT U116 ( .A1(MemOutputB3[26]), .A2(n3296), .A3(MemOutputB3[58]), 
        .A4(n3546), .A5(n69), .Y(n68) );
  AO22X1_RVT U117 ( .A1(MemOutputB3[90]), .A2(n3526), .A3(MemOutputB3[122]), 
        .A4(n3507), .Y(n69) );
  AO22X1_RVT U118 ( .A1(MemOutputB3[186]), .A2(n3258), .A3(MemOutputB3[154]), 
        .A4(n3283), .Y(n67) );
  AO22X1_RVT U119 ( .A1(MemOutputB3[218]), .A2(n3485), .A3(MemOutputB3[250]), 
        .A4(n3312), .Y(n66) );
  OR3X1_RVT U120 ( .A1(n70), .A2(n71), .A3(n72), .Y(ipB3[25]) );
  AO221X1_RVT U121 ( .A1(MemOutputB3[25]), .A2(n3308), .A3(MemOutputB3[57]), 
        .A4(n3546), .A5(n73), .Y(n72) );
  AO22X1_RVT U122 ( .A1(MemOutputB3[89]), .A2(n3526), .A3(MemOutputB3[121]), 
        .A4(n3507), .Y(n73) );
  AO22X1_RVT U123 ( .A1(MemOutputB3[185]), .A2(n3249), .A3(MemOutputB3[153]), 
        .A4(n454), .Y(n71) );
  AO22X1_RVT U124 ( .A1(MemOutputB3[217]), .A2(n3485), .A3(MemOutputB3[249]), 
        .A4(n3332), .Y(n70) );
  OR3X1_RVT U125 ( .A1(n74), .A2(n75), .A3(n76), .Y(ipB3[24]) );
  AO221X1_RVT U126 ( .A1(MemOutputB3[24]), .A2(n3305), .A3(MemOutputB3[56]), 
        .A4(n3546), .A5(n77), .Y(n76) );
  AO22X1_RVT U127 ( .A1(MemOutputB3[88]), .A2(n3526), .A3(MemOutputB3[120]), 
        .A4(n3507), .Y(n77) );
  AO22X1_RVT U128 ( .A1(MemOutputB3[184]), .A2(n3263), .A3(MemOutputB3[152]), 
        .A4(n3273), .Y(n75) );
  AO22X1_RVT U129 ( .A1(MemOutputB3[216]), .A2(n3485), .A3(MemOutputB3[248]), 
        .A4(n3332), .Y(n74) );
  OR3X1_RVT U130 ( .A1(n78), .A2(n79), .A3(n80), .Y(ipB3[23]) );
  AO221X1_RVT U131 ( .A1(MemOutputB3[23]), .A2(n3304), .A3(MemOutputB3[55]), 
        .A4(n3546), .A5(n81), .Y(n80) );
  AO22X1_RVT U132 ( .A1(MemOutputB3[87]), .A2(n3526), .A3(MemOutputB3[119]), 
        .A4(n3507), .Y(n81) );
  AO22X1_RVT U133 ( .A1(MemOutputB3[183]), .A2(n3262), .A3(MemOutputB3[151]), 
        .A4(n506), .Y(n79) );
  AO22X1_RVT U134 ( .A1(MemOutputB3[215]), .A2(n3485), .A3(MemOutputB3[247]), 
        .A4(n3333), .Y(n78) );
  OR3X1_RVT U135 ( .A1(n82), .A2(n83), .A3(n84), .Y(ipB3[22]) );
  AO221X1_RVT U136 ( .A1(MemOutputB3[22]), .A2(n3308), .A3(MemOutputB3[54]), 
        .A4(n3546), .A5(n85), .Y(n84) );
  AO22X1_RVT U137 ( .A1(MemOutputB3[86]), .A2(n3526), .A3(MemOutputB3[118]), 
        .A4(n3507), .Y(n85) );
  AO22X1_RVT U138 ( .A1(MemOutputB3[182]), .A2(n3265), .A3(MemOutputB3[150]), 
        .A4(n3286), .Y(n83) );
  AO22X1_RVT U139 ( .A1(MemOutputB3[214]), .A2(n3485), .A3(MemOutputB3[246]), 
        .A4(n3324), .Y(n82) );
  OR3X1_RVT U140 ( .A1(n86), .A2(n87), .A3(n88), .Y(ipB3[21]) );
  AO221X1_RVT U141 ( .A1(MemOutputB3[21]), .A2(n3304), .A3(MemOutputB3[53]), 
        .A4(n3546), .A5(n89), .Y(n88) );
  AO22X1_RVT U142 ( .A1(MemOutputB3[85]), .A2(n3526), .A3(MemOutputB3[117]), 
        .A4(n3507), .Y(n89) );
  AO22X1_RVT U143 ( .A1(MemOutputB3[181]), .A2(n3264), .A3(MemOutputB3[149]), 
        .A4(n3286), .Y(n87) );
  AO22X1_RVT U144 ( .A1(MemOutputB3[213]), .A2(n3485), .A3(MemOutputB3[245]), 
        .A4(n3332), .Y(n86) );
  OR3X1_RVT U145 ( .A1(n90), .A2(n91), .A3(n92), .Y(ipB3[20]) );
  AO221X1_RVT U146 ( .A1(MemOutputB3[20]), .A2(n3307), .A3(MemOutputB3[52]), 
        .A4(n3546), .A5(n93), .Y(n92) );
  AO22X1_RVT U147 ( .A1(MemOutputB3[84]), .A2(n3526), .A3(MemOutputB3[116]), 
        .A4(n3507), .Y(n93) );
  AO22X1_RVT U148 ( .A1(MemOutputB3[180]), .A2(n451), .A3(MemOutputB3[148]), 
        .A4(n454), .Y(n91) );
  AO22X1_RVT U149 ( .A1(MemOutputB3[212]), .A2(n3485), .A3(MemOutputB3[244]), 
        .A4(n3327), .Y(n90) );
  OR3X1_RVT U150 ( .A1(n94), .A2(n95), .A3(n96), .Y(ipB3[1]) );
  AO221X1_RVT U151 ( .A1(MemOutputB3[1]), .A2(n3307), .A3(MemOutputB3[33]), 
        .A4(n3546), .A5(n97), .Y(n96) );
  AO22X1_RVT U152 ( .A1(MemOutputB3[65]), .A2(n3526), .A3(MemOutputB3[97]), 
        .A4(n3507), .Y(n97) );
  AO22X1_RVT U153 ( .A1(MemOutputB3[161]), .A2(n3261), .A3(MemOutputB3[129]), 
        .A4(n3270), .Y(n95) );
  AO22X1_RVT U154 ( .A1(MemOutputB3[193]), .A2(n3485), .A3(MemOutputB3[225]), 
        .A4(n3329), .Y(n94) );
  OR3X1_RVT U155 ( .A1(n98), .A2(n99), .A3(n100), .Y(ipB3[19]) );
  AO221X1_RVT U156 ( .A1(MemOutputB3[19]), .A2(n3297), .A3(MemOutputB3[51]), 
        .A4(n3546), .A5(n101), .Y(n100) );
  AO22X1_RVT U157 ( .A1(MemOutputB3[83]), .A2(n3526), .A3(MemOutputB3[115]), 
        .A4(n3507), .Y(n101) );
  AO22X1_RVT U158 ( .A1(MemOutputB3[179]), .A2(n3253), .A3(MemOutputB3[147]), 
        .A4(n3279), .Y(n99) );
  AO22X1_RVT U159 ( .A1(MemOutputB3[211]), .A2(n3485), .A3(MemOutputB3[243]), 
        .A4(n3319), .Y(n98) );
  OR3X1_RVT U160 ( .A1(n102), .A2(n103), .A3(n104), .Y(ipB3[18]) );
  AO221X1_RVT U161 ( .A1(MemOutputB3[18]), .A2(n3302), .A3(MemOutputB3[50]), 
        .A4(n3546), .A5(n105), .Y(n104) );
  AO22X1_RVT U162 ( .A1(MemOutputB3[82]), .A2(n3526), .A3(MemOutputB3[114]), 
        .A4(n3507), .Y(n105) );
  AO22X1_RVT U163 ( .A1(MemOutputB3[178]), .A2(n3250), .A3(MemOutputB3[146]), 
        .A4(n3271), .Y(n103) );
  AO22X1_RVT U164 ( .A1(MemOutputB3[210]), .A2(n3485), .A3(MemOutputB3[242]), 
        .A4(n3316), .Y(n102) );
  OR3X1_RVT U165 ( .A1(n106), .A2(n107), .A3(n108), .Y(ipB3[17]) );
  AO221X1_RVT U166 ( .A1(MemOutputB3[17]), .A2(n3298), .A3(MemOutputB3[49]), 
        .A4(n3546), .A5(n109), .Y(n108) );
  AO22X1_RVT U167 ( .A1(MemOutputB3[81]), .A2(n3526), .A3(MemOutputB3[113]), 
        .A4(n3507), .Y(n109) );
  AO22X1_RVT U168 ( .A1(MemOutputB3[177]), .A2(n451), .A3(MemOutputB3[145]), 
        .A4(n506), .Y(n107) );
  AO22X1_RVT U169 ( .A1(MemOutputB3[209]), .A2(n3485), .A3(MemOutputB3[241]), 
        .A4(n3318), .Y(n106) );
  OR3X1_RVT U170 ( .A1(n110), .A2(n111), .A3(n112), .Y(ipB3[16]) );
  AO221X1_RVT U171 ( .A1(MemOutputB3[16]), .A2(n3298), .A3(MemOutputB3[48]), 
        .A4(n3547), .A5(n113), .Y(n112) );
  AO22X1_RVT U172 ( .A1(MemOutputB3[80]), .A2(n3527), .A3(MemOutputB3[112]), 
        .A4(n3508), .Y(n113) );
  AO22X1_RVT U173 ( .A1(MemOutputB3[176]), .A2(n3250), .A3(MemOutputB3[144]), 
        .A4(n3278), .Y(n111) );
  AO22X1_RVT U174 ( .A1(MemOutputB3[208]), .A2(n3486), .A3(MemOutputB3[240]), 
        .A4(n3316), .Y(n110) );
  OR3X1_RVT U175 ( .A1(n114), .A2(n115), .A3(n116), .Y(ipB3[15]) );
  AO221X1_RVT U176 ( .A1(MemOutputB3[15]), .A2(n3297), .A3(MemOutputB3[47]), 
        .A4(n3547), .A5(n117), .Y(n116) );
  AO22X1_RVT U177 ( .A1(MemOutputB3[79]), .A2(n3527), .A3(MemOutputB3[111]), 
        .A4(n3508), .Y(n117) );
  AO22X1_RVT U178 ( .A1(MemOutputB3[175]), .A2(n3265), .A3(MemOutputB3[143]), 
        .A4(n3288), .Y(n115) );
  AO22X1_RVT U179 ( .A1(MemOutputB3[207]), .A2(n3486), .A3(MemOutputB3[239]), 
        .A4(n3310), .Y(n114) );
  OR3X1_RVT U180 ( .A1(n118), .A2(n119), .A3(n120), .Y(ipB3[14]) );
  AO221X1_RVT U181 ( .A1(MemOutputB3[14]), .A2(n3297), .A3(MemOutputB3[46]), 
        .A4(n3547), .A5(n121), .Y(n120) );
  AO22X1_RVT U182 ( .A1(MemOutputB3[78]), .A2(n3527), .A3(MemOutputB3[110]), 
        .A4(n3508), .Y(n121) );
  AO22X1_RVT U183 ( .A1(MemOutputB3[174]), .A2(n3250), .A3(MemOutputB3[142]), 
        .A4(n3271), .Y(n119) );
  AO22X1_RVT U184 ( .A1(MemOutputB3[206]), .A2(n3486), .A3(MemOutputB3[238]), 
        .A4(n3313), .Y(n118) );
  OR3X1_RVT U185 ( .A1(n122), .A2(n123), .A3(n124), .Y(ipB3[13]) );
  AO221X1_RVT U186 ( .A1(MemOutputB3[13]), .A2(n3303), .A3(MemOutputB3[45]), 
        .A4(n3547), .A5(n125), .Y(n124) );
  AO22X1_RVT U187 ( .A1(MemOutputB3[77]), .A2(n3527), .A3(MemOutputB3[109]), 
        .A4(n3508), .Y(n125) );
  AO22X1_RVT U188 ( .A1(MemOutputB3[173]), .A2(n3249), .A3(MemOutputB3[141]), 
        .A4(n3270), .Y(n123) );
  OR3X1_RVT U190 ( .A1(n126), .A2(n127), .A3(n128), .Y(ipB3[12]) );
  AO221X1_RVT U191 ( .A1(MemOutputB3[12]), .A2(n3301), .A3(MemOutputB3[44]), 
        .A4(n3547), .A5(n129), .Y(n128) );
  AO22X1_RVT U192 ( .A1(MemOutputB3[76]), .A2(n3527), .A3(MemOutputB3[108]), 
        .A4(n3508), .Y(n129) );
  AO22X1_RVT U193 ( .A1(MemOutputB3[172]), .A2(n3254), .A3(MemOutputB3[140]), 
        .A4(n3273), .Y(n127) );
  AO22X1_RVT U194 ( .A1(MemOutputB3[204]), .A2(n3486), .A3(MemOutputB3[236]), 
        .A4(n3312), .Y(n126) );
  OR3X1_RVT U195 ( .A1(n130), .A2(n131), .A3(n132), .Y(ipB3[11]) );
  AO221X1_RVT U196 ( .A1(MemOutputB3[11]), .A2(n3298), .A3(MemOutputB3[43]), 
        .A4(n3547), .A5(n133), .Y(n132) );
  AO22X1_RVT U197 ( .A1(MemOutputB3[75]), .A2(n3527), .A3(MemOutputB3[107]), 
        .A4(n3508), .Y(n133) );
  AO22X1_RVT U198 ( .A1(MemOutputB3[171]), .A2(n3253), .A3(MemOutputB3[139]), 
        .A4(n506), .Y(n131) );
  AO22X1_RVT U199 ( .A1(MemOutputB3[203]), .A2(n3486), .A3(MemOutputB3[235]), 
        .A4(n3310), .Y(n130) );
  OR3X1_RVT U200 ( .A1(n134), .A2(n135), .A3(n136), .Y(ipB3[10]) );
  AO221X1_RVT U201 ( .A1(MemOutputB3[10]), .A2(n3298), .A3(MemOutputB3[42]), 
        .A4(n3547), .A5(n137), .Y(n136) );
  AO22X1_RVT U202 ( .A1(MemOutputB3[74]), .A2(n3527), .A3(MemOutputB3[106]), 
        .A4(n3508), .Y(n137) );
  AO22X1_RVT U203 ( .A1(MemOutputB3[170]), .A2(n3252), .A3(MemOutputB3[138]), 
        .A4(n506), .Y(n135) );
  AO22X1_RVT U204 ( .A1(MemOutputB3[202]), .A2(n3486), .A3(MemOutputB3[234]), 
        .A4(n3315), .Y(n134) );
  OR3X1_RVT U205 ( .A1(n138), .A2(n139), .A3(n140), .Y(ipB3[0]) );
  AO221X1_RVT U206 ( .A1(MemOutputB3[0]), .A2(n408), .A3(MemOutputB3[32]), 
        .A4(n3547), .A5(n141), .Y(n140) );
  AO22X1_RVT U207 ( .A1(MemOutputB3[64]), .A2(n3527), .A3(MemOutputB3[96]), 
        .A4(n3508), .Y(n141) );
  AO22X1_RVT U208 ( .A1(MemOutputB3[160]), .A2(n3262), .A3(MemOutputB3[128]), 
        .A4(n3283), .Y(n139) );
  AO22X1_RVT U209 ( .A1(MemOutputB3[192]), .A2(n3486), .A3(MemOutputB3[224]), 
        .A4(n3314), .Y(n138) );
  OR3X1_RVT U210 ( .A1(n142), .A2(n143), .A3(n144), .Y(ipB2[9]) );
  AO221X1_RVT U211 ( .A1(MemOutputB2[9]), .A2(n3296), .A3(MemOutputB2[41]), 
        .A4(n3547), .A5(n145), .Y(n144) );
  AO22X1_RVT U212 ( .A1(MemOutputB2[73]), .A2(n3527), .A3(MemOutputB2[105]), 
        .A4(n3508), .Y(n145) );
  AO22X1_RVT U213 ( .A1(MemOutputB2[169]), .A2(n3250), .A3(MemOutputB2[137]), 
        .A4(n3283), .Y(n143) );
  AO22X1_RVT U214 ( .A1(MemOutputB2[201]), .A2(n3486), .A3(MemOutputB2[233]), 
        .A4(n3315), .Y(n142) );
  OR3X1_RVT U215 ( .A1(n146), .A2(n147), .A3(n148), .Y(ipB2[8]) );
  AO221X1_RVT U216 ( .A1(MemOutputB2[8]), .A2(n3302), .A3(MemOutputB2[40]), 
        .A4(n3547), .A5(n149), .Y(n148) );
  AO22X1_RVT U217 ( .A1(MemOutputB2[72]), .A2(n3527), .A3(MemOutputB2[104]), 
        .A4(n3508), .Y(n149) );
  AO22X1_RVT U218 ( .A1(MemOutputB2[168]), .A2(n3258), .A3(MemOutputB2[136]), 
        .A4(n3281), .Y(n147) );
  AO22X1_RVT U219 ( .A1(MemOutputB2[200]), .A2(n3486), .A3(MemOutputB2[232]), 
        .A4(n3317), .Y(n146) );
  OR3X1_RVT U220 ( .A1(n150), .A2(n151), .A3(n152), .Y(ipB2[7]) );
  AO221X1_RVT U221 ( .A1(MemOutputB2[7]), .A2(n3297), .A3(MemOutputB2[39]), 
        .A4(n3547), .A5(n153), .Y(n152) );
  AO22X1_RVT U222 ( .A1(MemOutputB2[71]), .A2(n3527), .A3(MemOutputB2[103]), 
        .A4(n3508), .Y(n153) );
  AO22X1_RVT U223 ( .A1(MemOutputB2[167]), .A2(n3264), .A3(MemOutputB2[135]), 
        .A4(n3275), .Y(n151) );
  AO22X1_RVT U224 ( .A1(MemOutputB2[199]), .A2(n3486), .A3(MemOutputB2[231]), 
        .A4(n3312), .Y(n150) );
  OR3X1_RVT U225 ( .A1(n154), .A2(n155), .A3(n156), .Y(ipB2[6]) );
  AO221X1_RVT U226 ( .A1(MemOutputB2[6]), .A2(n3295), .A3(MemOutputB2[38]), 
        .A4(n3547), .A5(n157), .Y(n156) );
  AO22X1_RVT U227 ( .A1(MemOutputB2[70]), .A2(n3527), .A3(MemOutputB2[102]), 
        .A4(n3508), .Y(n157) );
  AO22X1_RVT U228 ( .A1(MemOutputB2[166]), .A2(n3264), .A3(MemOutputB2[134]), 
        .A4(n506), .Y(n155) );
  AO22X1_RVT U229 ( .A1(MemOutputB2[198]), .A2(n3486), .A3(MemOutputB2[230]), 
        .A4(n3312), .Y(n154) );
  OR3X1_RVT U230 ( .A1(n158), .A2(n159), .A3(n160), .Y(ipB2[5]) );
  AO221X1_RVT U231 ( .A1(MemOutputB2[5]), .A2(n3297), .A3(MemOutputB2[37]), 
        .A4(n3548), .A5(n161), .Y(n160) );
  AO22X1_RVT U232 ( .A1(MemOutputB2[69]), .A2(n3528), .A3(MemOutputB2[101]), 
        .A4(n3509), .Y(n161) );
  AO22X1_RVT U233 ( .A1(MemOutputB2[165]), .A2(n3249), .A3(MemOutputB2[133]), 
        .A4(n3283), .Y(n159) );
  AO22X1_RVT U234 ( .A1(MemOutputB2[197]), .A2(n3487), .A3(MemOutputB2[229]), 
        .A4(n3316), .Y(n158) );
  OR3X1_RVT U235 ( .A1(n162), .A2(n163), .A3(n164), .Y(ipB2[4]) );
  AO221X1_RVT U236 ( .A1(MemOutputB2[4]), .A2(n3307), .A3(MemOutputB2[36]), 
        .A4(n3548), .A5(n165), .Y(n164) );
  AO22X1_RVT U237 ( .A1(MemOutputB2[68]), .A2(n3528), .A3(MemOutputB2[100]), 
        .A4(n3509), .Y(n165) );
  AO22X1_RVT U238 ( .A1(MemOutputB2[164]), .A2(n3248), .A3(MemOutputB2[132]), 
        .A4(n3271), .Y(n163) );
  AO22X1_RVT U239 ( .A1(MemOutputB2[196]), .A2(n3487), .A3(MemOutputB2[228]), 
        .A4(n3310), .Y(n162) );
  OR3X1_RVT U240 ( .A1(n166), .A2(n167), .A3(n168), .Y(ipB2[3]) );
  AO221X1_RVT U241 ( .A1(MemOutputB2[3]), .A2(n3297), .A3(MemOutputB2[35]), 
        .A4(n3548), .A5(n169), .Y(n168) );
  AO22X1_RVT U242 ( .A1(MemOutputB2[67]), .A2(n3528), .A3(MemOutputB2[99]), 
        .A4(n3509), .Y(n169) );
  AO22X1_RVT U243 ( .A1(MemOutputB2[163]), .A2(n3248), .A3(MemOutputB2[131]), 
        .A4(n3277), .Y(n167) );
  AO22X1_RVT U244 ( .A1(MemOutputB2[195]), .A2(n3487), .A3(MemOutputB2[227]), 
        .A4(n3323), .Y(n166) );
  OR3X1_RVT U245 ( .A1(n170), .A2(n171), .A3(n172), .Y(ipB2[31]) );
  AO221X1_RVT U246 ( .A1(MemOutputB2[31]), .A2(n3302), .A3(MemOutputB2[63]), 
        .A4(n3548), .A5(n173), .Y(n172) );
  AO22X1_RVT U247 ( .A1(MemOutputB2[95]), .A2(n3528), .A3(MemOutputB2[127]), 
        .A4(n3509), .Y(n173) );
  AO22X1_RVT U248 ( .A1(MemOutputB2[191]), .A2(n514), .A3(MemOutputB2[159]), 
        .A4(n3276), .Y(n171) );
  AO22X1_RVT U249 ( .A1(MemOutputB2[223]), .A2(n3487), .A3(MemOutputB2[255]), 
        .A4(n3323), .Y(n170) );
  OR3X1_RVT U250 ( .A1(n174), .A2(n175), .A3(n176), .Y(ipB2[30]) );
  AO221X1_RVT U251 ( .A1(MemOutputB2[30]), .A2(n3299), .A3(MemOutputB2[62]), 
        .A4(n3548), .A5(n177), .Y(n176) );
  AO22X1_RVT U252 ( .A1(MemOutputB2[94]), .A2(n3528), .A3(MemOutputB2[126]), 
        .A4(n3509), .Y(n177) );
  AO22X1_RVT U254 ( .A1(MemOutputB2[222]), .A2(n3487), .A3(MemOutputB2[254]), 
        .A4(n3313), .Y(n174) );
  OR3X1_RVT U255 ( .A1(n178), .A2(n179), .A3(n180), .Y(ipB2[2]) );
  AO221X1_RVT U256 ( .A1(MemOutputB2[2]), .A2(n3298), .A3(MemOutputB2[34]), 
        .A4(n3548), .A5(n181), .Y(n180) );
  AO22X1_RVT U257 ( .A1(MemOutputB2[66]), .A2(n3528), .A3(MemOutputB2[98]), 
        .A4(n3509), .Y(n181) );
  AO22X1_RVT U258 ( .A1(MemOutputB2[162]), .A2(n514), .A3(MemOutputB2[130]), 
        .A4(n454), .Y(n179) );
  AO22X1_RVT U259 ( .A1(MemOutputB2[194]), .A2(n3487), .A3(MemOutputB2[226]), 
        .A4(n3322), .Y(n178) );
  OR3X1_RVT U260 ( .A1(n182), .A2(n183), .A3(n184), .Y(ipB2[29]) );
  AO221X1_RVT U261 ( .A1(MemOutputB2[29]), .A2(n3299), .A3(MemOutputB2[61]), 
        .A4(n3548), .A5(n185), .Y(n184) );
  AO22X1_RVT U262 ( .A1(MemOutputB2[93]), .A2(n3528), .A3(MemOutputB2[125]), 
        .A4(n3509), .Y(n185) );
  AO22X1_RVT U263 ( .A1(MemOutputB2[189]), .A2(n451), .A3(MemOutputB2[157]), 
        .A4(n3276), .Y(n183) );
  AO22X1_RVT U264 ( .A1(MemOutputB2[221]), .A2(n3487), .A3(MemOutputB2[253]), 
        .A4(n3325), .Y(n182) );
  OR3X1_RVT U265 ( .A1(n186), .A2(n187), .A3(n188), .Y(ipB2[28]) );
  AO221X1_RVT U266 ( .A1(MemOutputB2[28]), .A2(n3298), .A3(MemOutputB2[60]), 
        .A4(n3548), .A5(n189), .Y(n188) );
  AO22X1_RVT U267 ( .A1(MemOutputB2[92]), .A2(n3528), .A3(MemOutputB2[124]), 
        .A4(n3509), .Y(n189) );
  AO22X1_RVT U268 ( .A1(MemOutputB2[188]), .A2(n514), .A3(MemOutputB2[156]), 
        .A4(n3275), .Y(n187) );
  AO22X1_RVT U269 ( .A1(MemOutputB2[220]), .A2(n3487), .A3(MemOutputB2[252]), 
        .A4(n3318), .Y(n186) );
  OR3X1_RVT U270 ( .A1(n190), .A2(n191), .A3(n192), .Y(ipB2[27]) );
  AO221X1_RVT U271 ( .A1(MemOutputB2[27]), .A2(n3298), .A3(MemOutputB2[59]), 
        .A4(n3548), .A5(n193), .Y(n192) );
  AO22X1_RVT U272 ( .A1(MemOutputB2[91]), .A2(n3528), .A3(MemOutputB2[123]), 
        .A4(n3509), .Y(n193) );
  AO22X1_RVT U273 ( .A1(MemOutputB2[187]), .A2(n3249), .A3(MemOutputB2[155]), 
        .A4(n506), .Y(n191) );
  OR3X1_RVT U275 ( .A1(n194), .A2(n195), .A3(n196), .Y(ipB2[26]) );
  AO221X1_RVT U276 ( .A1(MemOutputB2[26]), .A2(n3298), .A3(MemOutputB2[58]), 
        .A4(n3548), .A5(n197), .Y(n196) );
  AO22X1_RVT U277 ( .A1(MemOutputB2[90]), .A2(n3528), .A3(MemOutputB2[122]), 
        .A4(n3509), .Y(n197) );
  AO22X1_RVT U278 ( .A1(MemOutputB2[186]), .A2(n3251), .A3(MemOutputB2[154]), 
        .A4(n3277), .Y(n195) );
  AO22X1_RVT U279 ( .A1(MemOutputB2[218]), .A2(n3487), .A3(MemOutputB2[250]), 
        .A4(n3324), .Y(n194) );
  OR3X1_RVT U280 ( .A1(n198), .A2(n199), .A3(n200), .Y(ipB2[25]) );
  AO221X1_RVT U281 ( .A1(MemOutputB2[25]), .A2(n3299), .A3(MemOutputB2[57]), 
        .A4(n3548), .A5(n201), .Y(n200) );
  AO22X1_RVT U282 ( .A1(MemOutputB2[89]), .A2(n3528), .A3(MemOutputB2[121]), 
        .A4(n3509), .Y(n201) );
  AO22X1_RVT U283 ( .A1(MemOutputB2[185]), .A2(n451), .A3(MemOutputB2[153]), 
        .A4(n506), .Y(n199) );
  AO22X1_RVT U284 ( .A1(MemOutputB2[217]), .A2(n3487), .A3(MemOutputB2[249]), 
        .A4(n3334), .Y(n198) );
  OR3X1_RVT U285 ( .A1(n202), .A2(n203), .A3(n204), .Y(ipB2[24]) );
  AO221X1_RVT U286 ( .A1(MemOutputB2[24]), .A2(n3298), .A3(MemOutputB2[56]), 
        .A4(n3548), .A5(n205), .Y(n204) );
  AO22X1_RVT U287 ( .A1(MemOutputB2[88]), .A2(n3528), .A3(MemOutputB2[120]), 
        .A4(n3509), .Y(n205) );
  AO22X1_RVT U288 ( .A1(MemOutputB2[184]), .A2(n3247), .A3(MemOutputB2[152]), 
        .A4(n3271), .Y(n203) );
  AO22X1_RVT U289 ( .A1(MemOutputB2[216]), .A2(n3487), .A3(MemOutputB2[248]), 
        .A4(n3324), .Y(n202) );
  OR3X1_RVT U290 ( .A1(n206), .A2(n207), .A3(n208), .Y(ipB2[23]) );
  AO221X1_RVT U291 ( .A1(MemOutputB2[23]), .A2(n3307), .A3(MemOutputB2[55]), 
        .A4(n3549), .A5(n209), .Y(n208) );
  AO22X1_RVT U292 ( .A1(MemOutputB2[87]), .A2(n3529), .A3(MemOutputB2[119]), 
        .A4(n3510), .Y(n209) );
  AO22X1_RVT U293 ( .A1(MemOutputB2[183]), .A2(n3249), .A3(MemOutputB2[151]), 
        .A4(n506), .Y(n207) );
  AO22X1_RVT U294 ( .A1(MemOutputB2[215]), .A2(n3488), .A3(MemOutputB2[247]), 
        .A4(n3334), .Y(n206) );
  OR3X1_RVT U295 ( .A1(n210), .A2(n211), .A3(n212), .Y(ipB2[22]) );
  AO221X1_RVT U296 ( .A1(MemOutputB2[22]), .A2(n3303), .A3(MemOutputB2[54]), 
        .A4(n3549), .A5(n213), .Y(n212) );
  AO22X1_RVT U297 ( .A1(MemOutputB2[86]), .A2(n3529), .A3(MemOutputB2[118]), 
        .A4(n3510), .Y(n213) );
  AO22X1_RVT U298 ( .A1(MemOutputB2[182]), .A2(n451), .A3(MemOutputB2[150]), 
        .A4(n3273), .Y(n211) );
  AO22X1_RVT U299 ( .A1(MemOutputB2[214]), .A2(n3488), .A3(MemOutputB2[246]), 
        .A4(n3330), .Y(n210) );
  OR3X1_RVT U300 ( .A1(n214), .A2(n215), .A3(n216), .Y(ipB2[21]) );
  AO221X1_RVT U301 ( .A1(MemOutputB2[21]), .A2(n3305), .A3(MemOutputB2[53]), 
        .A4(n3549), .A5(n217), .Y(n216) );
  AO22X1_RVT U302 ( .A1(MemOutputB2[85]), .A2(n3529), .A3(MemOutputB2[117]), 
        .A4(n3510), .Y(n217) );
  AO22X1_RVT U303 ( .A1(MemOutputB2[181]), .A2(n3247), .A3(MemOutputB2[149]), 
        .A4(n3282), .Y(n215) );
  AO22X1_RVT U304 ( .A1(MemOutputB2[213]), .A2(n3488), .A3(MemOutputB2[245]), 
        .A4(n3324), .Y(n214) );
  OR3X1_RVT U305 ( .A1(n218), .A2(n219), .A3(n220), .Y(ipB2[20]) );
  AO221X1_RVT U306 ( .A1(MemOutputB2[20]), .A2(n3307), .A3(MemOutputB2[52]), 
        .A4(n3549), .A5(n221), .Y(n220) );
  AO22X1_RVT U307 ( .A1(MemOutputB2[84]), .A2(n3529), .A3(MemOutputB2[116]), 
        .A4(n3510), .Y(n221) );
  AO22X1_RVT U308 ( .A1(MemOutputB2[180]), .A2(n3247), .A3(MemOutputB2[148]), 
        .A4(n3276), .Y(n219) );
  AO22X1_RVT U309 ( .A1(MemOutputB2[212]), .A2(n3488), .A3(MemOutputB2[244]), 
        .A4(n3327), .Y(n218) );
  OR3X1_RVT U310 ( .A1(n222), .A2(n223), .A3(n224), .Y(ipB2[1]) );
  AO221X1_RVT U311 ( .A1(MemOutputB2[1]), .A2(n3304), .A3(MemOutputB2[33]), 
        .A4(n3549), .A5(n225), .Y(n224) );
  AO22X1_RVT U312 ( .A1(MemOutputB2[65]), .A2(n3529), .A3(MemOutputB2[97]), 
        .A4(n3510), .Y(n225) );
  AO22X1_RVT U313 ( .A1(MemOutputB2[161]), .A2(n3262), .A3(MemOutputB2[129]), 
        .A4(n3281), .Y(n223) );
  AO22X1_RVT U314 ( .A1(MemOutputB2[193]), .A2(n3488), .A3(MemOutputB2[225]), 
        .A4(n3326), .Y(n222) );
  OR3X1_RVT U315 ( .A1(n226), .A2(n227), .A3(n228), .Y(ipB2[19]) );
  AO221X1_RVT U316 ( .A1(MemOutputB2[19]), .A2(n3297), .A3(MemOutputB2[51]), 
        .A4(n3549), .A5(n229), .Y(n228) );
  AO22X1_RVT U317 ( .A1(MemOutputB2[83]), .A2(n3529), .A3(MemOutputB2[115]), 
        .A4(n3510), .Y(n229) );
  AO22X1_RVT U318 ( .A1(MemOutputB2[179]), .A2(n3265), .A3(MemOutputB2[147]), 
        .A4(n454), .Y(n227) );
  AO22X1_RVT U319 ( .A1(MemOutputB2[211]), .A2(n3488), .A3(MemOutputB2[243]), 
        .A4(n3336), .Y(n226) );
  OR3X1_RVT U320 ( .A1(n230), .A2(n231), .A3(n232), .Y(ipB2[18]) );
  AO221X1_RVT U321 ( .A1(MemOutputB2[18]), .A2(n3304), .A3(MemOutputB2[50]), 
        .A4(n3549), .A5(n233), .Y(n232) );
  AO22X1_RVT U322 ( .A1(MemOutputB2[82]), .A2(n3529), .A3(MemOutputB2[114]), 
        .A4(n3510), .Y(n233) );
  AO22X1_RVT U323 ( .A1(MemOutputB2[178]), .A2(n3258), .A3(MemOutputB2[146]), 
        .A4(n3276), .Y(n231) );
  AO22X1_RVT U324 ( .A1(MemOutputB2[210]), .A2(n3488), .A3(MemOutputB2[242]), 
        .A4(n3327), .Y(n230) );
  OR3X1_RVT U325 ( .A1(n234), .A2(n235), .A3(n236), .Y(ipB2[17]) );
  AO221X1_RVT U326 ( .A1(MemOutputB2[17]), .A2(n3295), .A3(MemOutputB2[49]), 
        .A4(n3549), .A5(n237), .Y(n236) );
  AO22X1_RVT U327 ( .A1(MemOutputB2[81]), .A2(n3529), .A3(MemOutputB2[113]), 
        .A4(n3510), .Y(n237) );
  AO22X1_RVT U328 ( .A1(MemOutputB2[177]), .A2(n3247), .A3(MemOutputB2[145]), 
        .A4(n3277), .Y(n235) );
  AO22X1_RVT U329 ( .A1(MemOutputB2[209]), .A2(n3488), .A3(MemOutputB2[241]), 
        .A4(n3323), .Y(n234) );
  OR3X1_RVT U330 ( .A1(n238), .A2(n239), .A3(n240), .Y(ipB2[16]) );
  AO221X1_RVT U331 ( .A1(MemOutputB2[16]), .A2(n3304), .A3(MemOutputB2[48]), 
        .A4(n3549), .A5(n241), .Y(n240) );
  AO22X1_RVT U332 ( .A1(MemOutputB2[80]), .A2(n3529), .A3(MemOutputB2[112]), 
        .A4(n3510), .Y(n241) );
  AO22X1_RVT U333 ( .A1(MemOutputB2[176]), .A2(n3249), .A3(MemOutputB2[144]), 
        .A4(n3278), .Y(n239) );
  AO22X1_RVT U334 ( .A1(MemOutputB2[208]), .A2(n3488), .A3(MemOutputB2[240]), 
        .A4(n3326), .Y(n238) );
  OR3X1_RVT U335 ( .A1(n242), .A2(n243), .A3(n244), .Y(ipB2[15]) );
  AO221X1_RVT U336 ( .A1(MemOutputB2[15]), .A2(n3303), .A3(MemOutputB2[47]), 
        .A4(n3549), .A5(n245), .Y(n244) );
  AO22X1_RVT U337 ( .A1(MemOutputB2[79]), .A2(n3529), .A3(MemOutputB2[111]), 
        .A4(n3510), .Y(n245) );
  AO22X1_RVT U338 ( .A1(MemOutputB2[175]), .A2(n3254), .A3(MemOutputB2[143]), 
        .A4(n454), .Y(n243) );
  AO22X1_RVT U339 ( .A1(MemOutputB2[207]), .A2(n3488), .A3(MemOutputB2[239]), 
        .A4(n3319), .Y(n242) );
  OR3X1_RVT U340 ( .A1(n246), .A2(n247), .A3(n248), .Y(ipB2[14]) );
  AO221X1_RVT U341 ( .A1(MemOutputB2[14]), .A2(n3303), .A3(MemOutputB2[46]), 
        .A4(n3549), .A5(n249), .Y(n248) );
  AO22X1_RVT U342 ( .A1(MemOutputB2[78]), .A2(n3529), .A3(MemOutputB2[110]), 
        .A4(n3510), .Y(n249) );
  AO22X1_RVT U343 ( .A1(MemOutputB2[174]), .A2(n3253), .A3(MemOutputB2[142]), 
        .A4(n506), .Y(n247) );
  OR3X1_RVT U345 ( .A1(n250), .A2(n251), .A3(n252), .Y(ipB2[13]) );
  AO221X1_RVT U346 ( .A1(MemOutputB2[13]), .A2(n3307), .A3(MemOutputB2[45]), 
        .A4(n3549), .A5(n253), .Y(n252) );
  AO22X1_RVT U347 ( .A1(MemOutputB2[77]), .A2(n3529), .A3(MemOutputB2[109]), 
        .A4(n3510), .Y(n253) );
  AO22X1_RVT U348 ( .A1(MemOutputB2[173]), .A2(n3252), .A3(MemOutputB2[141]), 
        .A4(n3278), .Y(n251) );
  AO22X1_RVT U349 ( .A1(MemOutputB2[205]), .A2(n3488), .A3(MemOutputB2[237]), 
        .A4(n3319), .Y(n250) );
  OR3X1_RVT U350 ( .A1(n254), .A2(n255), .A3(n256), .Y(ipB2[12]) );
  AO221X1_RVT U351 ( .A1(MemOutputB2[12]), .A2(n3304), .A3(MemOutputB2[44]), 
        .A4(n3550), .A5(n257), .Y(n256) );
  AO22X1_RVT U352 ( .A1(MemOutputB2[76]), .A2(n3530), .A3(MemOutputB2[108]), 
        .A4(n3511), .Y(n257) );
  AO22X1_RVT U353 ( .A1(MemOutputB2[172]), .A2(n451), .A3(MemOutputB2[140]), 
        .A4(n3278), .Y(n255) );
  AO22X1_RVT U354 ( .A1(MemOutputB2[204]), .A2(n3489), .A3(MemOutputB2[236]), 
        .A4(n3319), .Y(n254) );
  OR3X1_RVT U355 ( .A1(n258), .A2(n259), .A3(n260), .Y(ipB2[11]) );
  AO221X1_RVT U356 ( .A1(MemOutputB2[11]), .A2(n3305), .A3(MemOutputB2[43]), 
        .A4(n3550), .A5(n261), .Y(n260) );
  AO22X1_RVT U357 ( .A1(MemOutputB2[75]), .A2(n3530), .A3(MemOutputB2[107]), 
        .A4(n3511), .Y(n261) );
  AO22X1_RVT U358 ( .A1(MemOutputB2[171]), .A2(n3257), .A3(MemOutputB2[139]), 
        .A4(n3277), .Y(n259) );
  AO22X1_RVT U359 ( .A1(MemOutputB2[203]), .A2(n3489), .A3(MemOutputB2[235]), 
        .A4(n3318), .Y(n258) );
  OR3X1_RVT U360 ( .A1(n262), .A2(n263), .A3(n264), .Y(ipB2[10]) );
  AO221X1_RVT U361 ( .A1(MemOutputB2[10]), .A2(n3303), .A3(MemOutputB2[42]), 
        .A4(n3550), .A5(n265), .Y(n264) );
  AO22X1_RVT U362 ( .A1(MemOutputB2[74]), .A2(n3530), .A3(MemOutputB2[106]), 
        .A4(n3511), .Y(n265) );
  AO22X1_RVT U363 ( .A1(MemOutputB2[170]), .A2(n3251), .A3(MemOutputB2[138]), 
        .A4(n3285), .Y(n263) );
  AO22X1_RVT U364 ( .A1(MemOutputB2[202]), .A2(n3489), .A3(MemOutputB2[234]), 
        .A4(n3315), .Y(n262) );
  OR3X1_RVT U365 ( .A1(n266), .A2(n267), .A3(n268), .Y(ipB2[0]) );
  AO221X1_RVT U366 ( .A1(MemOutputB2[0]), .A2(n3303), .A3(MemOutputB2[32]), 
        .A4(n3550), .A5(n269), .Y(n268) );
  AO22X1_RVT U367 ( .A1(MemOutputB2[64]), .A2(n3530), .A3(MemOutputB2[96]), 
        .A4(n3511), .Y(n269) );
  AO22X1_RVT U368 ( .A1(MemOutputB2[160]), .A2(n3262), .A3(MemOutputB2[128]), 
        .A4(n3283), .Y(n267) );
  AO22X1_RVT U369 ( .A1(MemOutputB2[192]), .A2(n3489), .A3(MemOutputB2[224]), 
        .A4(n3316), .Y(n266) );
  OR3X1_RVT U370 ( .A1(n270), .A2(n271), .A3(n272), .Y(ipB1[9]) );
  AO221X1_RVT U371 ( .A1(MemOutputB1[9]), .A2(n3297), .A3(MemOutputB1[41]), 
        .A4(n3550), .A5(n273), .Y(n272) );
  AO22X1_RVT U372 ( .A1(MemOutputB1[73]), .A2(n3530), .A3(MemOutputB1[105]), 
        .A4(n3511), .Y(n273) );
  AO22X1_RVT U373 ( .A1(MemOutputB1[169]), .A2(n3259), .A3(MemOutputB1[137]), 
        .A4(n3270), .Y(n271) );
  AO22X1_RVT U374 ( .A1(MemOutputB1[201]), .A2(n3489), .A3(MemOutputB1[233]), 
        .A4(n3316), .Y(n270) );
  OR3X1_RVT U375 ( .A1(n274), .A2(n275), .A3(n276), .Y(ipB1[8]) );
  AO221X1_RVT U376 ( .A1(MemOutputB1[8]), .A2(n3303), .A3(MemOutputB1[40]), 
        .A4(n3550), .A5(n277), .Y(n276) );
  AO22X1_RVT U377 ( .A1(MemOutputB1[72]), .A2(n3530), .A3(MemOutputB1[104]), 
        .A4(n3511), .Y(n277) );
  AO22X1_RVT U378 ( .A1(MemOutputB1[168]), .A2(n3257), .A3(MemOutputB1[136]), 
        .A4(n3272), .Y(n275) );
  AO22X1_RVT U379 ( .A1(MemOutputB1[200]), .A2(n3489), .A3(MemOutputB1[232]), 
        .A4(n3317), .Y(n274) );
  OR3X1_RVT U380 ( .A1(n278), .A2(n279), .A3(n280), .Y(ipB1[7]) );
  AO221X1_RVT U381 ( .A1(MemOutputB1[7]), .A2(n408), .A3(MemOutputB1[39]), 
        .A4(n3550), .A5(n281), .Y(n280) );
  AO22X1_RVT U382 ( .A1(MemOutputB1[71]), .A2(n3530), .A3(MemOutputB1[103]), 
        .A4(n3511), .Y(n281) );
  AO22X1_RVT U383 ( .A1(MemOutputB1[167]), .A2(n3262), .A3(MemOutputB1[135]), 
        .A4(n3272), .Y(n279) );
  AO22X1_RVT U384 ( .A1(MemOutputB1[199]), .A2(n3489), .A3(MemOutputB1[231]), 
        .A4(n3315), .Y(n278) );
  OR3X1_RVT U385 ( .A1(n282), .A2(n283), .A3(n284), .Y(ipB1[6]) );
  AO221X1_RVT U386 ( .A1(MemOutputB1[6]), .A2(n3301), .A3(MemOutputB1[38]), 
        .A4(n3550), .A5(n285), .Y(n284) );
  AO22X1_RVT U387 ( .A1(MemOutputB1[70]), .A2(n3530), .A3(MemOutputB1[102]), 
        .A4(n3511), .Y(n285) );
  AO22X1_RVT U388 ( .A1(MemOutputB1[166]), .A2(n451), .A3(MemOutputB1[134]), 
        .A4(n454), .Y(n283) );
  AO22X1_RVT U389 ( .A1(MemOutputB1[198]), .A2(n3489), .A3(MemOutputB1[230]), 
        .A4(n3312), .Y(n282) );
  OR3X1_RVT U390 ( .A1(n286), .A2(n287), .A3(n288), .Y(ipB1[5]) );
  AO221X1_RVT U391 ( .A1(MemOutputB1[5]), .A2(n3297), .A3(MemOutputB1[37]), 
        .A4(n3550), .A5(n289), .Y(n288) );
  AO22X1_RVT U392 ( .A1(MemOutputB1[69]), .A2(n3530), .A3(MemOutputB1[101]), 
        .A4(n3511), .Y(n289) );
  AO22X1_RVT U393 ( .A1(MemOutputB1[165]), .A2(n3261), .A3(MemOutputB1[133]), 
        .A4(n3278), .Y(n287) );
  AO22X1_RVT U394 ( .A1(MemOutputB1[197]), .A2(n3489), .A3(MemOutputB1[229]), 
        .A4(n3313), .Y(n286) );
  OR3X1_RVT U395 ( .A1(n290), .A2(n291), .A3(n292), .Y(ipB1[4]) );
  AO221X1_RVT U396 ( .A1(MemOutputB1[4]), .A2(n3307), .A3(MemOutputB1[36]), 
        .A4(n3550), .A5(n293), .Y(n292) );
  AO22X1_RVT U397 ( .A1(MemOutputB1[68]), .A2(n3530), .A3(MemOutputB1[100]), 
        .A4(n3511), .Y(n293) );
  AO22X1_RVT U398 ( .A1(MemOutputB1[164]), .A2(n3260), .A3(MemOutputB1[132]), 
        .A4(n506), .Y(n291) );
  AO22X1_RVT U399 ( .A1(MemOutputB1[196]), .A2(n3489), .A3(MemOutputB1[228]), 
        .A4(n3319), .Y(n290) );
  OR3X1_RVT U400 ( .A1(n294), .A2(n295), .A3(n296), .Y(ipB1[3]) );
  AO221X1_RVT U401 ( .A1(MemOutputB1[3]), .A2(n3297), .A3(MemOutputB1[35]), 
        .A4(n3550), .A5(n297), .Y(n296) );
  AO22X1_RVT U402 ( .A1(MemOutputB1[67]), .A2(n3530), .A3(MemOutputB1[99]), 
        .A4(n3511), .Y(n297) );
  AO22X1_RVT U403 ( .A1(MemOutputB1[163]), .A2(n3247), .A3(MemOutputB1[131]), 
        .A4(n3286), .Y(n295) );
  AO22X1_RVT U404 ( .A1(MemOutputB1[195]), .A2(n3489), .A3(MemOutputB1[227]), 
        .A4(n3314), .Y(n294) );
  OR3X1_RVT U405 ( .A1(n298), .A2(n299), .A3(n300), .Y(ipB1[31]) );
  AO221X1_RVT U406 ( .A1(MemOutputB1[31]), .A2(n3297), .A3(MemOutputB1[63]), 
        .A4(n3550), .A5(n301), .Y(n300) );
  AO22X1_RVT U407 ( .A1(MemOutputB1[95]), .A2(n3530), .A3(MemOutputB1[127]), 
        .A4(n3511), .Y(n301) );
  AO22X1_RVT U408 ( .A1(MemOutputB1[191]), .A2(n3264), .A3(MemOutputB1[159]), 
        .A4(n3272), .Y(n299) );
  AO22X1_RVT U409 ( .A1(MemOutputB1[223]), .A2(n3489), .A3(MemOutputB1[255]), 
        .A4(n3314), .Y(n298) );
  OR3X1_RVT U410 ( .A1(n302), .A2(n303), .A3(n304), .Y(ipB1[30]) );
  AO221X1_RVT U411 ( .A1(MemOutputB1[30]), .A2(n3296), .A3(MemOutputB1[62]), 
        .A4(n3551), .A5(n305), .Y(n304) );
  AO22X1_RVT U412 ( .A1(MemOutputB1[94]), .A2(n3531), .A3(MemOutputB1[126]), 
        .A4(n3512), .Y(n305) );
  AO22X1_RVT U413 ( .A1(MemOutputB1[190]), .A2(n3265), .A3(MemOutputB1[158]), 
        .A4(n3282), .Y(n303) );
  AO22X1_RVT U414 ( .A1(MemOutputB1[222]), .A2(n3490), .A3(MemOutputB1[254]), 
        .A4(n3314), .Y(n302) );
  OR3X1_RVT U415 ( .A1(n306), .A2(n307), .A3(n308), .Y(ipB1[2]) );
  AO221X1_RVT U416 ( .A1(MemOutputB1[2]), .A2(n3298), .A3(MemOutputB1[34]), 
        .A4(n3551), .A5(n309), .Y(n308) );
  AO22X1_RVT U417 ( .A1(MemOutputB1[66]), .A2(n3531), .A3(MemOutputB1[98]), 
        .A4(n3512), .Y(n309) );
  AO22X1_RVT U418 ( .A1(MemOutputB1[162]), .A2(n3249), .A3(MemOutputB1[130]), 
        .A4(n506), .Y(n307) );
  AO22X1_RVT U419 ( .A1(MemOutputB1[194]), .A2(n3490), .A3(MemOutputB1[226]), 
        .A4(n3313), .Y(n306) );
  OR3X1_RVT U420 ( .A1(n310), .A2(n311), .A3(n312), .Y(ipB1[29]) );
  AO221X1_RVT U421 ( .A1(MemOutputB1[29]), .A2(n3298), .A3(MemOutputB1[61]), 
        .A4(n3551), .A5(n313), .Y(n312) );
  AO22X1_RVT U422 ( .A1(MemOutputB1[93]), .A2(n3531), .A3(MemOutputB1[125]), 
        .A4(n3512), .Y(n313) );
  AO22X1_RVT U423 ( .A1(MemOutputB1[189]), .A2(n3261), .A3(MemOutputB1[157]), 
        .A4(n506), .Y(n311) );
  AO22X1_RVT U424 ( .A1(MemOutputB1[221]), .A2(n3490), .A3(MemOutputB1[253]), 
        .A4(n3310), .Y(n310) );
  OR3X1_RVT U425 ( .A1(n314), .A2(n315), .A3(n316), .Y(ipB1[28]) );
  AO221X1_RVT U426 ( .A1(MemOutputB1[28]), .A2(n3296), .A3(MemOutputB1[60]), 
        .A4(n3551), .A5(n317), .Y(n316) );
  AO22X1_RVT U427 ( .A1(MemOutputB1[92]), .A2(n3531), .A3(MemOutputB1[124]), 
        .A4(n3512), .Y(n317) );
  AO22X1_RVT U428 ( .A1(MemOutputB1[188]), .A2(n3260), .A3(MemOutputB1[156]), 
        .A4(n506), .Y(n315) );
  AO22X1_RVT U429 ( .A1(MemOutputB1[220]), .A2(n3490), .A3(MemOutputB1[252]), 
        .A4(n3318), .Y(n314) );
  OR3X1_RVT U430 ( .A1(n318), .A2(n319), .A3(n320), .Y(ipB1[27]) );
  AO221X1_RVT U431 ( .A1(MemOutputB1[27]), .A2(n3304), .A3(MemOutputB1[59]), 
        .A4(n3551), .A5(n321), .Y(n320) );
  AO22X1_RVT U432 ( .A1(MemOutputB1[91]), .A2(n3531), .A3(MemOutputB1[123]), 
        .A4(n3512), .Y(n321) );
  AO22X1_RVT U433 ( .A1(MemOutputB1[187]), .A2(n3264), .A3(MemOutputB1[155]), 
        .A4(n454), .Y(n319) );
  AO22X1_RVT U434 ( .A1(MemOutputB1[219]), .A2(n3490), .A3(MemOutputB1[251]), 
        .A4(n3313), .Y(n318) );
  OR3X1_RVT U435 ( .A1(n322), .A2(n323), .A3(n324), .Y(ipB1[26]) );
  AO221X1_RVT U436 ( .A1(MemOutputB1[26]), .A2(n3298), .A3(MemOutputB1[58]), 
        .A4(n3551), .A5(n325), .Y(n324) );
  AO22X1_RVT U437 ( .A1(MemOutputB1[90]), .A2(n3531), .A3(MemOutputB1[122]), 
        .A4(n3512), .Y(n325) );
  AO22X1_RVT U438 ( .A1(MemOutputB1[186]), .A2(n3250), .A3(MemOutputB1[154]), 
        .A4(n3279), .Y(n323) );
  AO22X1_RVT U439 ( .A1(MemOutputB1[218]), .A2(n3490), .A3(MemOutputB1[250]), 
        .A4(n3313), .Y(n322) );
  OR3X1_RVT U440 ( .A1(n326), .A2(n327), .A3(n328), .Y(ipB1[25]) );
  AO221X1_RVT U441 ( .A1(MemOutputB1[25]), .A2(n3291), .A3(MemOutputB1[57]), 
        .A4(n3551), .A5(n329), .Y(n328) );
  AO22X1_RVT U442 ( .A1(MemOutputB1[89]), .A2(n3531), .A3(MemOutputB1[121]), 
        .A4(n3512), .Y(n329) );
  AO22X1_RVT U443 ( .A1(MemOutputB1[185]), .A2(n3264), .A3(MemOutputB1[153]), 
        .A4(n3277), .Y(n327) );
  AO22X1_RVT U444 ( .A1(MemOutputB1[217]), .A2(n3490), .A3(MemOutputB1[249]), 
        .A4(n3326), .Y(n326) );
  OR3X1_RVT U445 ( .A1(n330), .A2(n331), .A3(n332), .Y(ipB1[24]) );
  AO221X1_RVT U446 ( .A1(MemOutputB1[24]), .A2(n3297), .A3(MemOutputB1[56]), 
        .A4(n3551), .A5(n333), .Y(n332) );
  AO22X1_RVT U447 ( .A1(MemOutputB1[88]), .A2(n3531), .A3(MemOutputB1[120]), 
        .A4(n3512), .Y(n333) );
  AO22X1_RVT U448 ( .A1(MemOutputB1[184]), .A2(n3262), .A3(MemOutputB1[152]), 
        .A4(n3285), .Y(n331) );
  AO22X1_RVT U449 ( .A1(MemOutputB1[216]), .A2(n3490), .A3(MemOutputB1[248]), 
        .A4(n3325), .Y(n330) );
  OR3X1_RVT U450 ( .A1(n334), .A2(n335), .A3(n336), .Y(ipB1[23]) );
  AO221X1_RVT U451 ( .A1(MemOutputB1[23]), .A2(n3297), .A3(MemOutputB1[55]), 
        .A4(n3551), .A5(n337), .Y(n336) );
  AO22X1_RVT U452 ( .A1(MemOutputB1[87]), .A2(n3531), .A3(MemOutputB1[119]), 
        .A4(n3512), .Y(n337) );
  AO22X1_RVT U453 ( .A1(MemOutputB1[183]), .A2(n451), .A3(MemOutputB1[151]), 
        .A4(n3275), .Y(n335) );
  AO22X1_RVT U454 ( .A1(MemOutputB1[215]), .A2(n3490), .A3(MemOutputB1[247]), 
        .A4(n3334), .Y(n334) );
  OR3X1_RVT U455 ( .A1(n338), .A2(n339), .A3(n340), .Y(ipB1[22]) );
  AO221X1_RVT U456 ( .A1(MemOutputB1[22]), .A2(n3302), .A3(MemOutputB1[54]), 
        .A4(n3551), .A5(n341), .Y(n340) );
  AO22X1_RVT U457 ( .A1(MemOutputB1[86]), .A2(n3531), .A3(MemOutputB1[118]), 
        .A4(n3512), .Y(n341) );
  AO22X1_RVT U458 ( .A1(MemOutputB1[182]), .A2(n3257), .A3(MemOutputB1[150]), 
        .A4(n506), .Y(n339) );
  AO22X1_RVT U459 ( .A1(MemOutputB1[214]), .A2(n3490), .A3(MemOutputB1[246]), 
        .A4(n3322), .Y(n338) );
  OR3X1_RVT U460 ( .A1(n342), .A2(n343), .A3(n344), .Y(ipB1[21]) );
  AO221X1_RVT U461 ( .A1(MemOutputB1[21]), .A2(n3291), .A3(MemOutputB1[53]), 
        .A4(n3551), .A5(n345), .Y(n344) );
  AO22X1_RVT U462 ( .A1(MemOutputB1[85]), .A2(n3531), .A3(MemOutputB1[117]), 
        .A4(n3512), .Y(n345) );
  AO22X1_RVT U463 ( .A1(MemOutputB1[181]), .A2(n3262), .A3(MemOutputB1[149]), 
        .A4(n3282), .Y(n343) );
  AO22X1_RVT U464 ( .A1(MemOutputB1[213]), .A2(n3490), .A3(MemOutputB1[245]), 
        .A4(n3322), .Y(n342) );
  OR3X1_RVT U465 ( .A1(n346), .A2(n347), .A3(n348), .Y(ipB1[20]) );
  AO221X1_RVT U466 ( .A1(MemOutputB1[20]), .A2(n3299), .A3(MemOutputB1[52]), 
        .A4(n3551), .A5(n349), .Y(n348) );
  AO22X1_RVT U467 ( .A1(MemOutputB1[84]), .A2(n3531), .A3(MemOutputB1[116]), 
        .A4(n3512), .Y(n349) );
  AO22X1_RVT U468 ( .A1(MemOutputB1[180]), .A2(n3248), .A3(MemOutputB1[148]), 
        .A4(n3270), .Y(n347) );
  AO22X1_RVT U469 ( .A1(MemOutputB1[212]), .A2(n3490), .A3(MemOutputB1[244]), 
        .A4(n3329), .Y(n346) );
  OR3X1_RVT U470 ( .A1(n350), .A2(n351), .A3(n352), .Y(ipB1[1]) );
  AO221X1_RVT U471 ( .A1(MemOutputB1[1]), .A2(n3297), .A3(MemOutputB1[33]), 
        .A4(n3552), .A5(n353), .Y(n352) );
  AO22X1_RVT U472 ( .A1(MemOutputB1[65]), .A2(n3527), .A3(MemOutputB1[97]), 
        .A4(n3513), .Y(n353) );
  AO22X1_RVT U473 ( .A1(MemOutputB1[161]), .A2(n3263), .A3(MemOutputB1[129]), 
        .A4(n3281), .Y(n351) );
  AO22X1_RVT U474 ( .A1(MemOutputB1[193]), .A2(n3491), .A3(MemOutputB1[225]), 
        .A4(n3336), .Y(n350) );
  OR3X1_RVT U475 ( .A1(n354), .A2(n355), .A3(n356), .Y(ipB1[19]) );
  AO221X1_RVT U476 ( .A1(MemOutputB1[19]), .A2(n3304), .A3(MemOutputB1[51]), 
        .A4(n3554), .A5(n357), .Y(n356) );
  AO22X1_RVT U477 ( .A1(MemOutputB1[83]), .A2(n3541), .A3(MemOutputB1[115]), 
        .A4(n3513), .Y(n357) );
  AO22X1_RVT U479 ( .A1(MemOutputB1[211]), .A2(n3491), .A3(MemOutputB1[243]), 
        .A4(n3333), .Y(n354) );
  OR3X1_RVT U480 ( .A1(n358), .A2(n359), .A3(n360), .Y(ipB1[18]) );
  AO221X1_RVT U481 ( .A1(MemOutputB1[18]), .A2(n3308), .A3(MemOutputB1[50]), 
        .A4(n3554), .A5(n361), .Y(n360) );
  AO22X1_RVT U482 ( .A1(MemOutputB1[82]), .A2(n519), .A3(MemOutputB1[114]), 
        .A4(n3513), .Y(n361) );
  AO22X1_RVT U483 ( .A1(MemOutputB1[178]), .A2(n3250), .A3(MemOutputB1[146]), 
        .A4(n3281), .Y(n359) );
  AO22X1_RVT U484 ( .A1(MemOutputB1[210]), .A2(n3491), .A3(MemOutputB1[242]), 
        .A4(n3327), .Y(n358) );
  OR3X1_RVT U485 ( .A1(n362), .A2(n363), .A3(n364), .Y(ipB1[17]) );
  AO221X1_RVT U486 ( .A1(MemOutputB1[17]), .A2(n3307), .A3(MemOutputB1[49]), 
        .A4(n3552), .A5(n365), .Y(n364) );
  AO22X1_RVT U487 ( .A1(MemOutputB1[81]), .A2(n3541), .A3(MemOutputB1[113]), 
        .A4(n3513), .Y(n365) );
  AO22X1_RVT U488 ( .A1(MemOutputB1[177]), .A2(n3257), .A3(MemOutputB1[145]), 
        .A4(n454), .Y(n363) );
  AO22X1_RVT U489 ( .A1(MemOutputB1[209]), .A2(n3491), .A3(MemOutputB1[241]), 
        .A4(n3318), .Y(n362) );
  OR3X1_RVT U490 ( .A1(n366), .A2(n367), .A3(n368), .Y(ipB1[16]) );
  AO221X1_RVT U491 ( .A1(MemOutputB1[16]), .A2(n3305), .A3(MemOutputB1[48]), 
        .A4(n3554), .A5(n369), .Y(n368) );
  AO22X1_RVT U492 ( .A1(MemOutputB1[80]), .A2(n507), .A3(MemOutputB1[112]), 
        .A4(n3513), .Y(n369) );
  AO22X1_RVT U493 ( .A1(MemOutputB1[176]), .A2(n3254), .A3(MemOutputB1[144]), 
        .A4(n3285), .Y(n367) );
  OR3X1_RVT U495 ( .A1(n370), .A2(n371), .A3(n372), .Y(ipB1[15]) );
  AO221X1_RVT U496 ( .A1(MemOutputB1[15]), .A2(n3297), .A3(MemOutputB1[47]), 
        .A4(n3552), .A5(n373), .Y(n372) );
  AO22X1_RVT U497 ( .A1(MemOutputB1[79]), .A2(n519), .A3(MemOutputB1[111]), 
        .A4(n3513), .Y(n373) );
  AO22X1_RVT U498 ( .A1(MemOutputB1[175]), .A2(n3253), .A3(MemOutputB1[143]), 
        .A4(n3286), .Y(n371) );
  AO22X1_RVT U499 ( .A1(MemOutputB1[207]), .A2(n3491), .A3(MemOutputB1[239]), 
        .A4(n3319), .Y(n370) );
  OR3X1_RVT U500 ( .A1(n374), .A2(n375), .A3(n376), .Y(ipB1[14]) );
  AO221X1_RVT U501 ( .A1(MemOutputB1[14]), .A2(n3307), .A3(MemOutputB1[46]), 
        .A4(n3554), .A5(n377), .Y(n376) );
  AO22X1_RVT U502 ( .A1(MemOutputB1[78]), .A2(n3541), .A3(MemOutputB1[110]), 
        .A4(n3513), .Y(n377) );
  AO22X1_RVT U503 ( .A1(MemOutputB1[174]), .A2(n3258), .A3(MemOutputB1[142]), 
        .A4(n3281), .Y(n375) );
  AO22X1_RVT U504 ( .A1(MemOutputB1[206]), .A2(n3491), .A3(MemOutputB1[238]), 
        .A4(n3320), .Y(n374) );
  OR3X1_RVT U505 ( .A1(n378), .A2(n379), .A3(n380), .Y(ipB1[13]) );
  AO221X1_RVT U506 ( .A1(MemOutputB1[13]), .A2(n3308), .A3(MemOutputB1[45]), 
        .A4(n3552), .A5(n381), .Y(n380) );
  AO22X1_RVT U507 ( .A1(MemOutputB1[77]), .A2(n507), .A3(MemOutputB1[109]), 
        .A4(n3513), .Y(n381) );
  AO22X1_RVT U508 ( .A1(MemOutputB1[173]), .A2(n451), .A3(MemOutputB1[141]), 
        .A4(n3279), .Y(n379) );
  AO22X1_RVT U509 ( .A1(MemOutputB1[205]), .A2(n3491), .A3(MemOutputB1[237]), 
        .A4(n3319), .Y(n378) );
  OR3X1_RVT U510 ( .A1(n382), .A2(n383), .A3(n384), .Y(ipB1[12]) );
  AO221X1_RVT U511 ( .A1(MemOutputB1[12]), .A2(n3298), .A3(MemOutputB1[44]), 
        .A4(n3554), .A5(n385), .Y(n384) );
  AO22X1_RVT U512 ( .A1(MemOutputB1[76]), .A2(n3538), .A3(MemOutputB1[108]), 
        .A4(n3513), .Y(n385) );
  AO22X1_RVT U513 ( .A1(MemOutputB1[172]), .A2(n3251), .A3(MemOutputB1[140]), 
        .A4(n3279), .Y(n383) );
  AO22X1_RVT U514 ( .A1(MemOutputB1[204]), .A2(n3491), .A3(MemOutputB1[236]), 
        .A4(n3317), .Y(n382) );
  OR3X1_RVT U515 ( .A1(n386), .A2(n387), .A3(n388), .Y(ipB1[11]) );
  AO221X1_RVT U516 ( .A1(MemOutputB1[11]), .A2(n3305), .A3(MemOutputB1[43]), 
        .A4(n3552), .A5(n389), .Y(n388) );
  AO22X1_RVT U517 ( .A1(MemOutputB1[75]), .A2(n507), .A3(MemOutputB1[107]), 
        .A4(n3513), .Y(n389) );
  AO22X1_RVT U518 ( .A1(MemOutputB1[171]), .A2(n3257), .A3(MemOutputB1[139]), 
        .A4(n3285), .Y(n387) );
  AO22X1_RVT U519 ( .A1(MemOutputB1[203]), .A2(n3491), .A3(MemOutputB1[235]), 
        .A4(n3314), .Y(n386) );
  OR3X1_RVT U520 ( .A1(n390), .A2(n391), .A3(n392), .Y(ipB1[10]) );
  AO221X1_RVT U521 ( .A1(MemOutputB1[10]), .A2(n3304), .A3(MemOutputB1[42]), 
        .A4(n3552), .A5(n393), .Y(n392) );
  AO22X1_RVT U522 ( .A1(MemOutputB1[74]), .A2(n3541), .A3(MemOutputB1[106]), 
        .A4(n3513), .Y(n393) );
  AO22X1_RVT U523 ( .A1(MemOutputB1[170]), .A2(n3265), .A3(MemOutputB1[138]), 
        .A4(n454), .Y(n391) );
  AO22X1_RVT U524 ( .A1(MemOutputB1[202]), .A2(n3491), .A3(MemOutputB1[234]), 
        .A4(n3317), .Y(n390) );
  OR3X1_RVT U525 ( .A1(n394), .A2(n395), .A3(n396), .Y(ipB1[0]) );
  AO221X1_RVT U526 ( .A1(MemOutputB1[0]), .A2(n3308), .A3(MemOutputB1[32]), 
        .A4(n3554), .A5(n397), .Y(n396) );
  AO22X1_RVT U527 ( .A1(MemOutputB1[64]), .A2(n519), .A3(MemOutputB1[96]), 
        .A4(n3513), .Y(n397) );
  AO22X1_RVT U528 ( .A1(MemOutputB1[160]), .A2(n3262), .A3(MemOutputB1[128]), 
        .A4(n3283), .Y(n395) );
  AO22X1_RVT U529 ( .A1(MemOutputB1[192]), .A2(n3491), .A3(MemOutputB1[224]), 
        .A4(n3315), .Y(n394) );
  AO22X1_RVT U532 ( .A1(MemOutputB0[73]), .A2(n3542), .A3(MemOutputB0[105]), 
        .A4(n935), .Y(n401) );
  AO22X1_RVT U537 ( .A1(MemOutputB0[72]), .A2(n3540), .A3(MemOutputB0[104]), 
        .A4(n934), .Y(n405) );
  AO221X1_RVT U546 ( .A1(MemOutputB0[6]), .A2(n3293), .A3(MemOutputB0[38]), 
        .A4(n10), .A5(n413), .Y(n412) );
  AO22X1_RVT U547 ( .A1(MemOutputB0[70]), .A2(n3540), .A3(MemOutputB0[102]), 
        .A4(n3522), .Y(n413) );
  AO22X1_RVT U548 ( .A1(MemOutputB0[166]), .A2(n3261), .A3(MemOutputB0[134]), 
        .A4(n3277), .Y(n411) );
  AO22X1_RVT U549 ( .A1(MemOutputB0[198]), .A2(n3492), .A3(MemOutputB0[230]), 
        .A4(n3327), .Y(n410) );
  OR3X1_RVT U550 ( .A1(n414), .A2(n415), .A3(n416), .Y(ipB0[5]) );
  AO221X1_RVT U551 ( .A1(MemOutputB0[5]), .A2(n456), .A3(MemOutputB0[37]), 
        .A4(n3564), .A5(n417), .Y(n416) );
  AO22X1_RVT U552 ( .A1(MemOutputB0[69]), .A2(n3542), .A3(MemOutputB0[101]), 
        .A4(n3515), .Y(n417) );
  AO22X1_RVT U553 ( .A1(MemOutputB0[165]), .A2(n3256), .A3(MemOutputB0[133]), 
        .A4(n3286), .Y(n415) );
  AO22X1_RVT U554 ( .A1(MemOutputB0[197]), .A2(n3492), .A3(MemOutputB0[229]), 
        .A4(n3323), .Y(n414) );
  OR3X1_RVT U560 ( .A1(n422), .A2(n423), .A3(n424), .Y(ipB0[3]) );
  AO221X1_RVT U561 ( .A1(MemOutputB0[3]), .A2(n3293), .A3(MemOutputB0[35]), 
        .A4(n3564), .A5(n425), .Y(n424) );
  AO22X1_RVT U562 ( .A1(MemOutputB0[67]), .A2(n3533), .A3(MemOutputB0[99]), 
        .A4(n934), .Y(n425) );
  AO22X1_RVT U563 ( .A1(MemOutputB0[163]), .A2(n3247), .A3(MemOutputB0[131]), 
        .A4(n3273), .Y(n423) );
  AO22X1_RVT U564 ( .A1(MemOutputB0[195]), .A2(n3492), .A3(MemOutputB0[227]), 
        .A4(n3315), .Y(n422) );
  OR3X1_RVT U565 ( .A1(n426), .A2(n427), .A3(n428), .Y(ipB0[31]) );
  AO221X1_RVT U566 ( .A1(MemOutputB0[31]), .A2(n3308), .A3(MemOutputB0[63]), 
        .A4(n3546), .A5(n429), .Y(n428) );
  AO22X1_RVT U568 ( .A1(MemOutputB0[191]), .A2(n3249), .A3(MemOutputB0[159]), 
        .A4(n3271), .Y(n427) );
  AO22X1_RVT U569 ( .A1(MemOutputB0[223]), .A2(n3492), .A3(MemOutputB0[255]), 
        .A4(n3326), .Y(n426) );
  AO221X1_RVT U571 ( .A1(MemOutputB0[30]), .A2(n3292), .A3(MemOutputB0[62]), 
        .A4(n3563), .A5(n433), .Y(n432) );
  AO22X1_RVT U573 ( .A1(MemOutputB0[190]), .A2(n3257), .A3(MemOutputB0[158]), 
        .A4(n3274), .Y(n431) );
  AO221X1_RVT U576 ( .A1(MemOutputB0[2]), .A2(n3295), .A3(MemOutputB0[34]), 
        .A4(n3562), .A5(n437), .Y(n436) );
  AO22X1_RVT U578 ( .A1(MemOutputB0[162]), .A2(n3259), .A3(MemOutputB0[130]), 
        .A4(n3275), .Y(n435) );
  AO22X1_RVT U579 ( .A1(MemOutputB0[194]), .A2(n3492), .A3(MemOutputB0[226]), 
        .A4(n3314), .Y(n434) );
  AO22X1_RVT U582 ( .A1(MemOutputB0[93]), .A2(n3241), .A3(MemOutputB0[125]), 
        .A4(n3523), .Y(n441) );
  AO22X1_RVT U587 ( .A1(MemOutputB0[92]), .A2(n3542), .A3(MemOutputB0[124]), 
        .A4(n3523), .Y(n445) );
  AO22X1_RVT U592 ( .A1(n3532), .A2(MemOutputB0[91]), .A3(MemOutputB0[123]), 
        .A4(n3514), .Y(n449) );
  AO22X1_RVT U597 ( .A1(n3241), .A2(MemOutputB0[90]), .A3(n3515), .A4(
        MemOutputB0[122]), .Y(n453) );
  AO22X1_RVT U602 ( .A1(n3533), .A2(MemOutputB0[89]), .A3(MemOutputB0[121]), 
        .A4(n3515), .Y(n457) );
  AO22X1_RVT U607 ( .A1(n3532), .A2(MemOutputB0[88]), .A3(n3514), .A4(
        MemOutputB0[120]), .Y(n461) );
  AO22X1_RVT U612 ( .A1(n3533), .A2(MemOutputB0[87]), .A3(MemOutputB0[119]), 
        .A4(n3236), .Y(n465) );
  AO22X1_RVT U617 ( .A1(n3532), .A2(MemOutputB0[86]), .A3(MemOutputB0[118]), 
        .A4(n508), .Y(n469) );
  AO22X1_RVT U622 ( .A1(n3532), .A2(MemOutputB0[85]), .A3(MemOutputB0[117]), 
        .A4(n508), .Y(n473) );
  AO22X1_RVT U627 ( .A1(n3532), .A2(MemOutputB0[84]), .A3(n3514), .A4(
        MemOutputB0[116]), .Y(n477) );
  OR3X1_RVT U630 ( .A1(n478), .A2(n479), .A3(n480), .Y(ipB0[1]) );
  AO221X1_RVT U631 ( .A1(MemOutputB0[1]), .A2(n456), .A3(MemOutputB0[33]), 
        .A4(n3562), .A5(n481), .Y(n480) );
  AO22X1_RVT U632 ( .A1(MemOutputB0[65]), .A2(n3542), .A3(MemOutputB0[97]), 
        .A4(n3515), .Y(n481) );
  AO22X1_RVT U633 ( .A1(MemOutputB0[161]), .A2(n3250), .A3(MemOutputB0[129]), 
        .A4(n3288), .Y(n479) );
  AO22X1_RVT U634 ( .A1(MemOutputB0[193]), .A2(n3505), .A3(MemOutputB0[225]), 
        .A4(n3318), .Y(n478) );
  AO22X1_RVT U637 ( .A1(MemOutputB0[83]), .A2(n3241), .A3(n3515), .A4(
        MemOutputB0[115]), .Y(n485) );
  AO22X1_RVT U642 ( .A1(MemOutputB0[82]), .A2(n3241), .A3(MemOutputB0[114]), 
        .A4(n3236), .Y(n489) );
  AO22X1_RVT U647 ( .A1(MemOutputB0[81]), .A2(n3241), .A3(MemOutputB0[113]), 
        .A4(n508), .Y(n493) );
  AO22X1_RVT U652 ( .A1(MemOutputB0[80]), .A2(n3533), .A3(MemOutputB0[112]), 
        .A4(n3515), .Y(n497) );
  AO22X1_RVT U672 ( .A1(MemOutputB0[76]), .A2(n3533), .A3(MemOutputB0[108]), 
        .A4(n3515), .Y(n513) );
  AO22X1_RVT U677 ( .A1(MemOutputB0[75]), .A2(n3241), .A3(MemOutputB0[107]), 
        .A4(n508), .Y(n517) );
  AO22X1_RVT U687 ( .A1(MemOutputB0[64]), .A2(n15), .A3(MemOutputB0[96]), .A4(
        n3522), .Y(n525) );
  OR3X1_RVT U690 ( .A1(n526), .A2(n527), .A3(n528), .Y(ipA3[9]) );
  AO221X1_RVT U691 ( .A1(MemOutputA3[9]), .A2(n3298), .A3(MemOutputA3[41]), 
        .A4(n3554), .A5(n529), .Y(n528) );
  AO22X1_RVT U692 ( .A1(MemOutputA3[73]), .A2(n519), .A3(MemOutputA3[105]), 
        .A4(n3518), .Y(n529) );
  AO22X1_RVT U693 ( .A1(MemOutputA3[169]), .A2(n3257), .A3(MemOutputA3[137]), 
        .A4(n3271), .Y(n527) );
  AO22X1_RVT U694 ( .A1(MemOutputA3[201]), .A2(n3486), .A3(MemOutputA3[233]), 
        .A4(n3327), .Y(n526) );
  OR3X1_RVT U695 ( .A1(n530), .A2(n531), .A3(n532), .Y(ipA3[8]) );
  AO221X1_RVT U696 ( .A1(MemOutputA3[8]), .A2(n3296), .A3(MemOutputA3[40]), 
        .A4(n3554), .A5(n533), .Y(n532) );
  AO22X1_RVT U697 ( .A1(MemOutputA3[72]), .A2(n519), .A3(MemOutputA3[104]), 
        .A4(n3512), .Y(n533) );
  AO22X1_RVT U698 ( .A1(MemOutputA3[168]), .A2(n3254), .A3(MemOutputA3[136]), 
        .A4(n3285), .Y(n531) );
  AO22X1_RVT U699 ( .A1(MemOutputA3[200]), .A2(n3494), .A3(MemOutputA3[232]), 
        .A4(n3329), .Y(n530) );
  OR3X1_RVT U700 ( .A1(n534), .A2(n535), .A3(n536), .Y(ipA3[7]) );
  AO221X1_RVT U701 ( .A1(MemOutputA3[7]), .A2(n3301), .A3(MemOutputA3[39]), 
        .A4(n3552), .A5(n537), .Y(n536) );
  AO22X1_RVT U703 ( .A1(MemOutputA3[167]), .A2(n3251), .A3(MemOutputA3[135]), 
        .A4(n3275), .Y(n535) );
  AO22X1_RVT U704 ( .A1(MemOutputA3[199]), .A2(n3490), .A3(MemOutputA3[231]), 
        .A4(n3336), .Y(n534) );
  OR3X1_RVT U705 ( .A1(n538), .A2(n539), .A3(n540), .Y(ipA3[6]) );
  AO221X1_RVT U706 ( .A1(MemOutputA3[6]), .A2(n3295), .A3(MemOutputA3[38]), 
        .A4(n3552), .A5(n541), .Y(n540) );
  AO22X1_RVT U708 ( .A1(MemOutputA3[166]), .A2(n3252), .A3(MemOutputA3[134]), 
        .A4(n3276), .Y(n539) );
  AO22X1_RVT U709 ( .A1(MemOutputA3[198]), .A2(n3489), .A3(MemOutputA3[230]), 
        .A4(n3330), .Y(n538) );
  OR3X1_RVT U710 ( .A1(n542), .A2(n543), .A3(n544), .Y(ipA3[5]) );
  AO221X1_RVT U711 ( .A1(MemOutputA3[5]), .A2(n3297), .A3(MemOutputA3[37]), 
        .A4(n3552), .A5(n545), .Y(n544) );
  AO22X1_RVT U712 ( .A1(MemOutputA3[69]), .A2(n507), .A3(MemOutputA3[101]), 
        .A4(n3516), .Y(n545) );
  AO22X1_RVT U713 ( .A1(MemOutputA3[165]), .A2(n514), .A3(MemOutputA3[133]), 
        .A4(n3288), .Y(n543) );
  AO22X1_RVT U714 ( .A1(MemOutputA3[197]), .A2(n3493), .A3(MemOutputA3[229]), 
        .A4(n3322), .Y(n542) );
  OR3X1_RVT U715 ( .A1(n546), .A2(n547), .A3(n548), .Y(ipA3[4]) );
  AO221X1_RVT U716 ( .A1(MemOutputA3[4]), .A2(n3295), .A3(MemOutputA3[36]), 
        .A4(n3554), .A5(n549), .Y(n548) );
  AO22X1_RVT U717 ( .A1(MemOutputA3[68]), .A2(n3539), .A3(MemOutputA3[100]), 
        .A4(n3516), .Y(n549) );
  AO22X1_RVT U718 ( .A1(MemOutputA3[164]), .A2(n3249), .A3(MemOutputA3[132]), 
        .A4(n3283), .Y(n547) );
  AO22X1_RVT U719 ( .A1(MemOutputA3[196]), .A2(n3493), .A3(MemOutputA3[228]), 
        .A4(n3322), .Y(n546) );
  OR3X1_RVT U720 ( .A1(n550), .A2(n551), .A3(n552), .Y(ipA3[3]) );
  AO221X1_RVT U721 ( .A1(MemOutputA3[3]), .A2(n3304), .A3(MemOutputA3[35]), 
        .A4(n3552), .A5(n553), .Y(n552) );
  AO22X1_RVT U722 ( .A1(MemOutputA3[67]), .A2(n507), .A3(MemOutputA3[99]), 
        .A4(n3516), .Y(n553) );
  AO22X1_RVT U723 ( .A1(MemOutputA3[163]), .A2(n3247), .A3(MemOutputA3[131]), 
        .A4(n3277), .Y(n551) );
  AO22X1_RVT U724 ( .A1(MemOutputA3[195]), .A2(n3493), .A3(MemOutputA3[227]), 
        .A4(n3315), .Y(n550) );
  OR3X1_RVT U725 ( .A1(n554), .A2(n555), .A3(n556), .Y(ipA3[31]) );
  AO221X1_RVT U726 ( .A1(MemOutputA3[31]), .A2(n3297), .A3(MemOutputA3[63]), 
        .A4(n3554), .A5(n557), .Y(n556) );
  AO22X1_RVT U727 ( .A1(MemOutputA3[95]), .A2(n3541), .A3(MemOutputA3[127]), 
        .A4(n3516), .Y(n557) );
  AO22X1_RVT U728 ( .A1(MemOutputA3[191]), .A2(n3247), .A3(MemOutputA3[159]), 
        .A4(n3272), .Y(n555) );
  AO22X1_RVT U729 ( .A1(MemOutputA3[223]), .A2(n3493), .A3(MemOutputA3[255]), 
        .A4(n3336), .Y(n554) );
  OR3X1_RVT U730 ( .A1(n558), .A2(n559), .A3(n560), .Y(ipA3[30]) );
  AO221X1_RVT U731 ( .A1(MemOutputA3[30]), .A2(n3299), .A3(MemOutputA3[62]), 
        .A4(n3554), .A5(n561), .Y(n560) );
  AO22X1_RVT U732 ( .A1(MemOutputA3[94]), .A2(n519), .A3(MemOutputA3[126]), 
        .A4(n3516), .Y(n561) );
  AO22X1_RVT U734 ( .A1(MemOutputA3[222]), .A2(n3493), .A3(MemOutputA3[254]), 
        .A4(n3320), .Y(n558) );
  OR3X1_RVT U735 ( .A1(n562), .A2(n563), .A3(n564), .Y(ipA3[2]) );
  AO221X1_RVT U736 ( .A1(MemOutputA3[2]), .A2(n3298), .A3(MemOutputA3[34]), 
        .A4(n3552), .A5(n565), .Y(n564) );
  AO22X1_RVT U737 ( .A1(MemOutputA3[66]), .A2(n519), .A3(MemOutputA3[98]), 
        .A4(n3516), .Y(n565) );
  AO22X1_RVT U738 ( .A1(MemOutputA3[162]), .A2(n3248), .A3(MemOutputA3[130]), 
        .A4(n3270), .Y(n563) );
  OR3X1_RVT U740 ( .A1(n566), .A2(n567), .A3(n568), .Y(ipA3[29]) );
  AO221X1_RVT U741 ( .A1(MemOutputA3[29]), .A2(n3299), .A3(MemOutputA3[61]), 
        .A4(n3554), .A5(n569), .Y(n568) );
  AO22X1_RVT U742 ( .A1(MemOutputA3[93]), .A2(n3541), .A3(MemOutputA3[125]), 
        .A4(n3516), .Y(n569) );
  AO22X1_RVT U743 ( .A1(MemOutputA3[189]), .A2(n3249), .A3(MemOutputA3[157]), 
        .A4(n454), .Y(n567) );
  AO22X1_RVT U744 ( .A1(MemOutputA3[221]), .A2(n3493), .A3(MemOutputA3[253]), 
        .A4(n3319), .Y(n566) );
  OR3X1_RVT U745 ( .A1(n570), .A2(n571), .A3(n572), .Y(ipA3[28]) );
  AO221X1_RVT U746 ( .A1(MemOutputA3[28]), .A2(n3298), .A3(MemOutputA3[60]), 
        .A4(n3552), .A5(n573), .Y(n572) );
  AO22X1_RVT U747 ( .A1(MemOutputA3[92]), .A2(n3538), .A3(MemOutputA3[124]), 
        .A4(n3516), .Y(n573) );
  AO22X1_RVT U748 ( .A1(MemOutputA3[188]), .A2(n3258), .A3(MemOutputA3[156]), 
        .A4(n3277), .Y(n571) );
  AO22X1_RVT U749 ( .A1(MemOutputA3[220]), .A2(n3493), .A3(MemOutputA3[252]), 
        .A4(n3319), .Y(n570) );
  OR3X1_RVT U750 ( .A1(n574), .A2(n575), .A3(n576), .Y(ipA3[27]) );
  AO221X1_RVT U751 ( .A1(MemOutputA3[27]), .A2(n3298), .A3(MemOutputA3[59]), 
        .A4(n3554), .A5(n577), .Y(n576) );
  AO22X1_RVT U752 ( .A1(MemOutputA3[91]), .A2(n3539), .A3(MemOutputA3[123]), 
        .A4(n3516), .Y(n577) );
  AO22X1_RVT U753 ( .A1(MemOutputA3[187]), .A2(n3259), .A3(MemOutputA3[155]), 
        .A4(n3281), .Y(n575) );
  AO22X1_RVT U754 ( .A1(MemOutputA3[219]), .A2(n3493), .A3(MemOutputA3[251]), 
        .A4(n3319), .Y(n574) );
  OR3X1_RVT U755 ( .A1(n578), .A2(n579), .A3(n580), .Y(ipA3[26]) );
  AO221X1_RVT U756 ( .A1(MemOutputA3[26]), .A2(n3297), .A3(MemOutputA3[58]), 
        .A4(n3552), .A5(n581), .Y(n580) );
  AO22X1_RVT U757 ( .A1(MemOutputA3[90]), .A2(n3539), .A3(MemOutputA3[122]), 
        .A4(n3516), .Y(n581) );
  AO22X1_RVT U758 ( .A1(MemOutputA3[186]), .A2(n514), .A3(MemOutputA3[154]), 
        .A4(n3276), .Y(n579) );
  AO22X1_RVT U759 ( .A1(MemOutputA3[218]), .A2(n3493), .A3(MemOutputA3[250]), 
        .A4(n3315), .Y(n578) );
  OR3X1_RVT U760 ( .A1(n582), .A2(n583), .A3(n584), .Y(ipA3[25]) );
  AO221X1_RVT U761 ( .A1(MemOutputA3[25]), .A2(n3291), .A3(MemOutputA3[57]), 
        .A4(n3554), .A5(n585), .Y(n584) );
  AO22X1_RVT U762 ( .A1(MemOutputA3[89]), .A2(n3528), .A3(MemOutputA3[121]), 
        .A4(n3516), .Y(n585) );
  AO22X1_RVT U763 ( .A1(MemOutputA3[185]), .A2(n451), .A3(MemOutputA3[153]), 
        .A4(n3272), .Y(n583) );
  AO22X1_RVT U764 ( .A1(MemOutputA3[217]), .A2(n3493), .A3(MemOutputA3[249]), 
        .A4(n3317), .Y(n582) );
  OR3X1_RVT U765 ( .A1(n586), .A2(n587), .A3(n588), .Y(ipA3[24]) );
  AO221X1_RVT U766 ( .A1(MemOutputA3[24]), .A2(n3303), .A3(MemOutputA3[56]), 
        .A4(n3552), .A5(n589), .Y(n588) );
  AO22X1_RVT U767 ( .A1(MemOutputA3[88]), .A2(n519), .A3(MemOutputA3[120]), 
        .A4(n3516), .Y(n589) );
  AO22X1_RVT U768 ( .A1(MemOutputA3[184]), .A2(n451), .A3(MemOutputA3[152]), 
        .A4(n3271), .Y(n587) );
  AO22X1_RVT U769 ( .A1(MemOutputA3[216]), .A2(n3493), .A3(MemOutputA3[248]), 
        .A4(n3330), .Y(n586) );
  OR3X1_RVT U770 ( .A1(n590), .A2(n591), .A3(n592), .Y(ipA3[23]) );
  AO221X1_RVT U771 ( .A1(MemOutputA3[23]), .A2(n3297), .A3(MemOutputA3[55]), 
        .A4(n3555), .A5(n593), .Y(n592) );
  AO22X1_RVT U772 ( .A1(MemOutputA3[87]), .A2(n3534), .A3(MemOutputA3[119]), 
        .A4(n3517), .Y(n593) );
  AO22X1_RVT U773 ( .A1(MemOutputA3[183]), .A2(n3261), .A3(MemOutputA3[151]), 
        .A4(n506), .Y(n591) );
  AO22X1_RVT U774 ( .A1(MemOutputA3[215]), .A2(n3494), .A3(MemOutputA3[247]), 
        .A4(n3326), .Y(n590) );
  OR3X1_RVT U775 ( .A1(n594), .A2(n595), .A3(n596), .Y(ipA3[22]) );
  AO221X1_RVT U776 ( .A1(MemOutputA3[22]), .A2(n3302), .A3(MemOutputA3[54]), 
        .A4(n3555), .A5(n597), .Y(n596) );
  AO22X1_RVT U777 ( .A1(MemOutputA3[86]), .A2(n3534), .A3(MemOutputA3[118]), 
        .A4(n3517), .Y(n597) );
  AO22X1_RVT U778 ( .A1(MemOutputA3[182]), .A2(n3260), .A3(MemOutputA3[150]), 
        .A4(n506), .Y(n595) );
  AO22X1_RVT U779 ( .A1(MemOutputA3[214]), .A2(n3494), .A3(MemOutputA3[246]), 
        .A4(n3326), .Y(n594) );
  OR3X1_RVT U780 ( .A1(n598), .A2(n599), .A3(n600), .Y(ipA3[21]) );
  AO221X1_RVT U781 ( .A1(MemOutputA3[21]), .A2(n3295), .A3(MemOutputA3[53]), 
        .A4(n3555), .A5(n601), .Y(n600) );
  AO22X1_RVT U782 ( .A1(MemOutputA3[85]), .A2(n3534), .A3(MemOutputA3[117]), 
        .A4(n3517), .Y(n601) );
  AO22X1_RVT U783 ( .A1(MemOutputA3[181]), .A2(n3257), .A3(MemOutputA3[149]), 
        .A4(n506), .Y(n599) );
  AO22X1_RVT U784 ( .A1(MemOutputA3[213]), .A2(n3494), .A3(MemOutputA3[245]), 
        .A4(n3329), .Y(n598) );
  OR3X1_RVT U785 ( .A1(n602), .A2(n603), .A3(n604), .Y(ipA3[20]) );
  AO221X1_RVT U786 ( .A1(MemOutputA3[20]), .A2(n3298), .A3(MemOutputA3[52]), 
        .A4(n3555), .A5(n605), .Y(n604) );
  AO22X1_RVT U787 ( .A1(MemOutputA3[84]), .A2(n3534), .A3(MemOutputA3[116]), 
        .A4(n3517), .Y(n605) );
  AO22X1_RVT U788 ( .A1(MemOutputA3[180]), .A2(n3252), .A3(MemOutputA3[148]), 
        .A4(n3288), .Y(n603) );
  AO22X1_RVT U789 ( .A1(MemOutputA3[212]), .A2(n3494), .A3(MemOutputA3[244]), 
        .A4(n3325), .Y(n602) );
  OR3X1_RVT U790 ( .A1(n606), .A2(n607), .A3(n608), .Y(ipA3[1]) );
  AO221X1_RVT U791 ( .A1(MemOutputA3[1]), .A2(n3296), .A3(MemOutputA3[33]), 
        .A4(n3555), .A5(n609), .Y(n608) );
  AO22X1_RVT U792 ( .A1(MemOutputA3[65]), .A2(n3534), .A3(MemOutputA3[97]), 
        .A4(n3517), .Y(n609) );
  AO22X1_RVT U793 ( .A1(MemOutputA3[161]), .A2(n3259), .A3(MemOutputA3[129]), 
        .A4(n3271), .Y(n607) );
  AO22X1_RVT U794 ( .A1(MemOutputA3[193]), .A2(n3494), .A3(MemOutputA3[225]), 
        .A4(n3332), .Y(n606) );
  OR3X1_RVT U795 ( .A1(n610), .A2(n611), .A3(n612), .Y(ipA3[19]) );
  AO221X1_RVT U796 ( .A1(MemOutputA3[19]), .A2(n3297), .A3(MemOutputA3[51]), 
        .A4(n3555), .A5(n613), .Y(n612) );
  AO22X1_RVT U797 ( .A1(MemOutputA3[83]), .A2(n3534), .A3(MemOutputA3[115]), 
        .A4(n3517), .Y(n613) );
  AO22X1_RVT U798 ( .A1(MemOutputA3[179]), .A2(n3262), .A3(MemOutputA3[147]), 
        .A4(n3288), .Y(n611) );
  AO22X1_RVT U799 ( .A1(MemOutputA3[211]), .A2(n3494), .A3(MemOutputA3[243]), 
        .A4(n3322), .Y(n610) );
  OR3X1_RVT U800 ( .A1(n614), .A2(n615), .A3(n616), .Y(ipA3[18]) );
  AO221X1_RVT U801 ( .A1(MemOutputA3[18]), .A2(n3298), .A3(MemOutputA3[50]), 
        .A4(n3555), .A5(n617), .Y(n616) );
  AO22X1_RVT U802 ( .A1(MemOutputA3[82]), .A2(n3534), .A3(MemOutputA3[114]), 
        .A4(n3517), .Y(n617) );
  AO22X1_RVT U803 ( .A1(MemOutputA3[178]), .A2(n3256), .A3(MemOutputA3[146]), 
        .A4(n3286), .Y(n615) );
  AO22X1_RVT U804 ( .A1(MemOutputA3[210]), .A2(n3494), .A3(MemOutputA3[242]), 
        .A4(n3322), .Y(n614) );
  OR3X1_RVT U805 ( .A1(n618), .A2(n619), .A3(n620), .Y(ipA3[17]) );
  AO221X1_RVT U806 ( .A1(MemOutputA3[17]), .A2(n3303), .A3(MemOutputA3[49]), 
        .A4(n3555), .A5(n621), .Y(n620) );
  AO22X1_RVT U807 ( .A1(MemOutputA3[81]), .A2(n3534), .A3(MemOutputA3[113]), 
        .A4(n3517), .Y(n621) );
  AO22X1_RVT U808 ( .A1(MemOutputA3[177]), .A2(n3251), .A3(MemOutputA3[145]), 
        .A4(n3288), .Y(n619) );
  AO22X1_RVT U809 ( .A1(MemOutputA3[209]), .A2(n3494), .A3(MemOutputA3[241]), 
        .A4(n3325), .Y(n618) );
  OR3X1_RVT U810 ( .A1(n622), .A2(n623), .A3(n624), .Y(ipA3[16]) );
  AO221X1_RVT U811 ( .A1(MemOutputA3[16]), .A2(n3297), .A3(MemOutputA3[48]), 
        .A4(n3555), .A5(n625), .Y(n624) );
  AO22X1_RVT U812 ( .A1(MemOutputA3[80]), .A2(n3534), .A3(MemOutputA3[112]), 
        .A4(n3517), .Y(n625) );
  AO22X1_RVT U813 ( .A1(MemOutputA3[176]), .A2(n3257), .A3(MemOutputA3[144]), 
        .A4(n3271), .Y(n623) );
  AO22X1_RVT U814 ( .A1(MemOutputA3[208]), .A2(n3494), .A3(MemOutputA3[240]), 
        .A4(n3322), .Y(n622) );
  OR3X1_RVT U815 ( .A1(n626), .A2(n627), .A3(n628), .Y(ipA3[15]) );
  AO221X1_RVT U816 ( .A1(MemOutputA3[15]), .A2(n3297), .A3(MemOutputA3[47]), 
        .A4(n3555), .A5(n629), .Y(n628) );
  AO22X1_RVT U817 ( .A1(MemOutputA3[79]), .A2(n3534), .A3(MemOutputA3[111]), 
        .A4(n3517), .Y(n629) );
  AO22X1_RVT U818 ( .A1(MemOutputA3[175]), .A2(n3263), .A3(MemOutputA3[143]), 
        .A4(n452), .Y(n627) );
  AO22X1_RVT U819 ( .A1(MemOutputA3[207]), .A2(n3494), .A3(MemOutputA3[239]), 
        .A4(n3327), .Y(n626) );
  OR3X1_RVT U820 ( .A1(n630), .A2(n631), .A3(n632), .Y(ipA3[14]) );
  AO221X1_RVT U821 ( .A1(MemOutputA3[14]), .A2(n3298), .A3(MemOutputA3[46]), 
        .A4(n3555), .A5(n633), .Y(n632) );
  AO22X1_RVT U822 ( .A1(MemOutputA3[78]), .A2(n3534), .A3(MemOutputA3[110]), 
        .A4(n3517), .Y(n633) );
  AO22X1_RVT U823 ( .A1(MemOutputA3[174]), .A2(n3249), .A3(MemOutputA3[142]), 
        .A4(n3277), .Y(n631) );
  AO22X1_RVT U824 ( .A1(MemOutputA3[206]), .A2(n3494), .A3(MemOutputA3[238]), 
        .A4(n3323), .Y(n630) );
  OR3X1_RVT U825 ( .A1(n634), .A2(n635), .A3(n636), .Y(ipA3[13]) );
  AO221X1_RVT U826 ( .A1(MemOutputA3[13]), .A2(n3298), .A3(MemOutputA3[45]), 
        .A4(n3555), .A5(n637), .Y(n636) );
  AO22X1_RVT U827 ( .A1(MemOutputA3[77]), .A2(n3534), .A3(MemOutputA3[109]), 
        .A4(n3517), .Y(n637) );
  AO22X1_RVT U828 ( .A1(MemOutputA3[173]), .A2(n3252), .A3(MemOutputA3[141]), 
        .A4(n3288), .Y(n635) );
  AO22X1_RVT U829 ( .A1(MemOutputA3[205]), .A2(n3494), .A3(MemOutputA3[237]), 
        .A4(n3329), .Y(n634) );
  OR3X1_RVT U830 ( .A1(n638), .A2(n639), .A3(n640), .Y(ipA3[12]) );
  AO221X1_RVT U831 ( .A1(MemOutputA3[12]), .A2(n3299), .A3(MemOutputA3[44]), 
        .A4(n3556), .A5(n641), .Y(n640) );
  AO22X1_RVT U832 ( .A1(MemOutputA3[76]), .A2(n3535), .A3(MemOutputA3[108]), 
        .A4(n3518), .Y(n641) );
  AO22X1_RVT U833 ( .A1(MemOutputA3[172]), .A2(n3264), .A3(MemOutputA3[140]), 
        .A4(n3278), .Y(n639) );
  AO22X1_RVT U834 ( .A1(MemOutputA3[204]), .A2(n3495), .A3(MemOutputA3[236]), 
        .A4(n3319), .Y(n638) );
  OR3X1_RVT U835 ( .A1(n642), .A2(n643), .A3(n644), .Y(ipA3[11]) );
  AO221X1_RVT U836 ( .A1(MemOutputA3[11]), .A2(n3298), .A3(MemOutputA3[43]), 
        .A4(n3556), .A5(n645), .Y(n644) );
  AO22X1_RVT U837 ( .A1(MemOutputA3[75]), .A2(n3535), .A3(MemOutputA3[107]), 
        .A4(n3518), .Y(n645) );
  AO22X1_RVT U838 ( .A1(MemOutputA3[171]), .A2(n3254), .A3(MemOutputA3[139]), 
        .A4(n3278), .Y(n643) );
  OR3X1_RVT U840 ( .A1(n646), .A2(n647), .A3(n648), .Y(ipA3[10]) );
  AO221X1_RVT U841 ( .A1(MemOutputA3[10]), .A2(n3299), .A3(MemOutputA3[42]), 
        .A4(n3556), .A5(n649), .Y(n648) );
  AO22X1_RVT U842 ( .A1(MemOutputA3[74]), .A2(n3535), .A3(MemOutputA3[106]), 
        .A4(n3518), .Y(n649) );
  AO22X1_RVT U843 ( .A1(MemOutputA3[170]), .A2(n3253), .A3(MemOutputA3[138]), 
        .A4(n3278), .Y(n647) );
  AO22X1_RVT U844 ( .A1(MemOutputA3[202]), .A2(n3495), .A3(MemOutputA3[234]), 
        .A4(n3320), .Y(n646) );
  OR3X1_RVT U845 ( .A1(n650), .A2(n651), .A3(n652), .Y(ipA3[0]) );
  AO221X1_RVT U846 ( .A1(MemOutputA3[0]), .A2(n3298), .A3(MemOutputA3[32]), 
        .A4(n3556), .A5(n653), .Y(n652) );
  AO22X1_RVT U847 ( .A1(MemOutputA3[64]), .A2(n3535), .A3(MemOutputA3[96]), 
        .A4(n3518), .Y(n653) );
  AO22X1_RVT U848 ( .A1(MemOutputA3[160]), .A2(n3250), .A3(MemOutputA3[128]), 
        .A4(n3279), .Y(n651) );
  AO22X1_RVT U849 ( .A1(MemOutputA3[192]), .A2(n3495), .A3(MemOutputA3[224]), 
        .A4(n3319), .Y(n650) );
  OR3X1_RVT U850 ( .A1(n654), .A2(n655), .A3(n656), .Y(ipA2[9]) );
  AO221X1_RVT U851 ( .A1(MemOutputA2[9]), .A2(n3298), .A3(MemOutputA2[41]), 
        .A4(n3556), .A5(n657), .Y(n656) );
  AO22X1_RVT U852 ( .A1(MemOutputA2[73]), .A2(n3535), .A3(MemOutputA2[105]), 
        .A4(n3518), .Y(n657) );
  AO22X1_RVT U853 ( .A1(MemOutputA2[169]), .A2(n451), .A3(MemOutputA2[137]), 
        .A4(n506), .Y(n655) );
  AO22X1_RVT U854 ( .A1(MemOutputA2[201]), .A2(n3495), .A3(MemOutputA2[233]), 
        .A4(n3320), .Y(n654) );
  OR3X1_RVT U855 ( .A1(n658), .A2(n659), .A3(n660), .Y(ipA2[8]) );
  AO221X1_RVT U856 ( .A1(MemOutputA2[8]), .A2(n3297), .A3(MemOutputA2[40]), 
        .A4(n3556), .A5(n661), .Y(n660) );
  AO22X1_RVT U857 ( .A1(MemOutputA2[72]), .A2(n3535), .A3(MemOutputA2[104]), 
        .A4(n3518), .Y(n661) );
  AO22X1_RVT U858 ( .A1(MemOutputA2[168]), .A2(n514), .A3(MemOutputA2[136]), 
        .A4(n454), .Y(n659) );
  AO22X1_RVT U859 ( .A1(MemOutputA2[200]), .A2(n3495), .A3(MemOutputA2[232]), 
        .A4(n3314), .Y(n658) );
  OR3X1_RVT U860 ( .A1(n662), .A2(n663), .A3(n664), .Y(ipA2[7]) );
  AO221X1_RVT U861 ( .A1(MemOutputA2[7]), .A2(n3304), .A3(MemOutputA2[39]), 
        .A4(n3556), .A5(n665), .Y(n664) );
  AO22X1_RVT U862 ( .A1(MemOutputA2[71]), .A2(n3535), .A3(MemOutputA2[103]), 
        .A4(n3518), .Y(n665) );
  AO22X1_RVT U863 ( .A1(MemOutputA2[167]), .A2(n3249), .A3(MemOutputA2[135]), 
        .A4(n3285), .Y(n663) );
  AO22X1_RVT U864 ( .A1(MemOutputA2[199]), .A2(n3495), .A3(MemOutputA2[231]), 
        .A4(n3333), .Y(n662) );
  OR3X1_RVT U865 ( .A1(n666), .A2(n667), .A3(n668), .Y(ipA2[6]) );
  AO221X1_RVT U866 ( .A1(MemOutputA2[6]), .A2(n3303), .A3(MemOutputA2[38]), 
        .A4(n3556), .A5(n669), .Y(n668) );
  AO22X1_RVT U867 ( .A1(MemOutputA2[70]), .A2(n3535), .A3(MemOutputA2[102]), 
        .A4(n3518), .Y(n669) );
  AO22X1_RVT U868 ( .A1(MemOutputA2[166]), .A2(n3258), .A3(MemOutputA2[134]), 
        .A4(n454), .Y(n667) );
  AO22X1_RVT U869 ( .A1(MemOutputA2[198]), .A2(n3495), .A3(MemOutputA2[230]), 
        .A4(n3336), .Y(n666) );
  OR3X1_RVT U870 ( .A1(n670), .A2(n671), .A3(n672), .Y(ipA2[5]) );
  AO221X1_RVT U871 ( .A1(MemOutputA2[5]), .A2(n3304), .A3(MemOutputA2[37]), 
        .A4(n3556), .A5(n673), .Y(n672) );
  AO22X1_RVT U872 ( .A1(MemOutputA2[69]), .A2(n3535), .A3(MemOutputA2[101]), 
        .A4(n3518), .Y(n673) );
  AO22X1_RVT U873 ( .A1(MemOutputA2[165]), .A2(n3249), .A3(MemOutputA2[133]), 
        .A4(n3279), .Y(n671) );
  AO22X1_RVT U874 ( .A1(MemOutputA2[197]), .A2(n3495), .A3(MemOutputA2[229]), 
        .A4(n3329), .Y(n670) );
  OR3X1_RVT U875 ( .A1(n674), .A2(n675), .A3(n676), .Y(ipA2[4]) );
  AO221X1_RVT U876 ( .A1(MemOutputA2[4]), .A2(n3302), .A3(MemOutputA2[36]), 
        .A4(n3556), .A5(n677), .Y(n676) );
  AO22X1_RVT U877 ( .A1(MemOutputA2[68]), .A2(n3535), .A3(MemOutputA2[100]), 
        .A4(n3518), .Y(n677) );
  AO22X1_RVT U878 ( .A1(MemOutputA2[164]), .A2(n3262), .A3(MemOutputA2[132]), 
        .A4(n506), .Y(n675) );
  AO22X1_RVT U879 ( .A1(MemOutputA2[196]), .A2(n3495), .A3(MemOutputA2[228]), 
        .A4(n3329), .Y(n674) );
  OR3X1_RVT U880 ( .A1(n678), .A2(n679), .A3(n680), .Y(ipA2[3]) );
  AO221X1_RVT U881 ( .A1(MemOutputA2[3]), .A2(n3298), .A3(MemOutputA2[35]), 
        .A4(n3556), .A5(n681), .Y(n680) );
  AO22X1_RVT U882 ( .A1(MemOutputA2[67]), .A2(n3535), .A3(MemOutputA2[99]), 
        .A4(n3518), .Y(n681) );
  AO22X1_RVT U883 ( .A1(MemOutputA2[163]), .A2(n451), .A3(MemOutputA2[131]), 
        .A4(n3283), .Y(n679) );
  AO22X1_RVT U884 ( .A1(MemOutputA2[195]), .A2(n3495), .A3(MemOutputA2[227]), 
        .A4(n3327), .Y(n678) );
  OR3X1_RVT U885 ( .A1(n682), .A2(n683), .A3(n684), .Y(ipA2[31]) );
  AO221X1_RVT U886 ( .A1(MemOutputA2[31]), .A2(n3297), .A3(MemOutputA2[63]), 
        .A4(n3556), .A5(n685), .Y(n684) );
  AO22X1_RVT U887 ( .A1(MemOutputA2[95]), .A2(n3535), .A3(MemOutputA2[127]), 
        .A4(n3518), .Y(n685) );
  AO22X1_RVT U888 ( .A1(MemOutputA2[191]), .A2(n3262), .A3(MemOutputA2[159]), 
        .A4(n454), .Y(n683) );
  AO22X1_RVT U889 ( .A1(MemOutputA2[223]), .A2(n3495), .A3(MemOutputA2[255]), 
        .A4(n3330), .Y(n682) );
  OR3X1_RVT U890 ( .A1(n686), .A2(n687), .A3(n688), .Y(ipA2[30]) );
  AO221X1_RVT U891 ( .A1(MemOutputA2[30]), .A2(n3307), .A3(MemOutputA2[62]), 
        .A4(n3557), .A5(n689), .Y(n688) );
  AO22X1_RVT U892 ( .A1(MemOutputA2[94]), .A2(n3536), .A3(MemOutputA2[126]), 
        .A4(n3510), .Y(n689) );
  AO22X1_RVT U893 ( .A1(MemOutputA2[190]), .A2(n3260), .A3(MemOutputA2[158]), 
        .A4(n3279), .Y(n687) );
  AO22X1_RVT U894 ( .A1(MemOutputA2[222]), .A2(n3496), .A3(MemOutputA2[254]), 
        .A4(n3320), .Y(n686) );
  OR3X1_RVT U895 ( .A1(n690), .A2(n691), .A3(n692), .Y(ipA2[2]) );
  AO221X1_RVT U896 ( .A1(MemOutputA2[2]), .A2(n3305), .A3(MemOutputA2[34]), 
        .A4(n3557), .A5(n693), .Y(n692) );
  AO22X1_RVT U897 ( .A1(MemOutputA2[66]), .A2(n3536), .A3(MemOutputA2[98]), 
        .A4(n3512), .Y(n693) );
  AO22X1_RVT U898 ( .A1(MemOutputA2[162]), .A2(n3259), .A3(MemOutputA2[130]), 
        .A4(n506), .Y(n691) );
  AO22X1_RVT U899 ( .A1(MemOutputA2[194]), .A2(n3496), .A3(MemOutputA2[226]), 
        .A4(n3318), .Y(n690) );
  OR3X1_RVT U900 ( .A1(n694), .A2(n695), .A3(n696), .Y(ipA2[29]) );
  AO221X1_RVT U901 ( .A1(MemOutputA2[29]), .A2(n3308), .A3(MemOutputA2[61]), 
        .A4(n3557), .A5(n697), .Y(n696) );
  AO22X1_RVT U902 ( .A1(MemOutputA2[93]), .A2(n3536), .A3(MemOutputA2[125]), 
        .A4(n3508), .Y(n697) );
  AO22X1_RVT U903 ( .A1(MemOutputA2[189]), .A2(n3250), .A3(MemOutputA2[157]), 
        .A4(n3283), .Y(n695) );
  AO22X1_RVT U904 ( .A1(MemOutputA2[221]), .A2(n3496), .A3(MemOutputA2[253]), 
        .A4(n3318), .Y(n694) );
  OR3X1_RVT U905 ( .A1(n698), .A2(n699), .A3(n700), .Y(ipA2[28]) );
  AO221X1_RVT U906 ( .A1(MemOutputA2[28]), .A2(n3303), .A3(MemOutputA2[60]), 
        .A4(n3557), .A5(n701), .Y(n700) );
  AO22X1_RVT U907 ( .A1(MemOutputA2[92]), .A2(n3536), .A3(MemOutputA2[124]), 
        .A4(n3518), .Y(n701) );
  AO22X1_RVT U908 ( .A1(MemOutputA2[188]), .A2(n3259), .A3(MemOutputA2[156]), 
        .A4(n3271), .Y(n699) );
  AO22X1_RVT U909 ( .A1(MemOutputA2[220]), .A2(n3496), .A3(MemOutputA2[252]), 
        .A4(n3317), .Y(n698) );
  OR3X1_RVT U910 ( .A1(n702), .A2(n703), .A3(n704), .Y(ipA2[27]) );
  AO221X1_RVT U911 ( .A1(MemOutputA2[27]), .A2(n3308), .A3(MemOutputA2[59]), 
        .A4(n3557), .A5(n705), .Y(n704) );
  AO22X1_RVT U912 ( .A1(MemOutputA2[91]), .A2(n3536), .A3(MemOutputA2[123]), 
        .A4(n3508), .Y(n705) );
  AO22X1_RVT U913 ( .A1(MemOutputA2[187]), .A2(n3262), .A3(MemOutputA2[155]), 
        .A4(n3286), .Y(n703) );
  AO22X1_RVT U914 ( .A1(MemOutputA2[219]), .A2(n3496), .A3(MemOutputA2[251]), 
        .A4(n3316), .Y(n702) );
  OR3X1_RVT U915 ( .A1(n706), .A2(n707), .A3(n708), .Y(ipA2[26]) );
  AO221X1_RVT U916 ( .A1(MemOutputA2[26]), .A2(n3304), .A3(MemOutputA2[58]), 
        .A4(n3557), .A5(n709), .Y(n708) );
  AO22X1_RVT U917 ( .A1(MemOutputA2[90]), .A2(n3536), .A3(MemOutputA2[122]), 
        .A4(n3509), .Y(n709) );
  AO22X1_RVT U918 ( .A1(MemOutputA2[186]), .A2(n451), .A3(MemOutputA2[154]), 
        .A4(n3275), .Y(n707) );
  AO22X1_RVT U919 ( .A1(MemOutputA2[218]), .A2(n3496), .A3(MemOutputA2[250]), 
        .A4(n3316), .Y(n706) );
  OR3X1_RVT U920 ( .A1(n710), .A2(n711), .A3(n712), .Y(ipA2[25]) );
  AO221X1_RVT U921 ( .A1(MemOutputA2[25]), .A2(n3298), .A3(MemOutputA2[57]), 
        .A4(n3557), .A5(n713), .Y(n712) );
  AO22X1_RVT U922 ( .A1(MemOutputA2[89]), .A2(n3536), .A3(MemOutputA2[121]), 
        .A4(n3509), .Y(n713) );
  AO22X1_RVT U923 ( .A1(MemOutputA2[185]), .A2(n3263), .A3(MemOutputA2[153]), 
        .A4(n506), .Y(n711) );
  AO22X1_RVT U924 ( .A1(MemOutputA2[217]), .A2(n3496), .A3(MemOutputA2[249]), 
        .A4(n3315), .Y(n710) );
  OR3X1_RVT U925 ( .A1(n714), .A2(n715), .A3(n716), .Y(ipA2[24]) );
  AO221X1_RVT U926 ( .A1(MemOutputA2[24]), .A2(n3297), .A3(MemOutputA2[56]), 
        .A4(n3557), .A5(n717), .Y(n716) );
  AO22X1_RVT U927 ( .A1(MemOutputA2[88]), .A2(n3536), .A3(MemOutputA2[120]), 
        .A4(n3508), .Y(n717) );
  AO22X1_RVT U928 ( .A1(MemOutputA2[184]), .A2(n3263), .A3(MemOutputA2[152]), 
        .A4(n3271), .Y(n715) );
  AO22X1_RVT U929 ( .A1(MemOutputA2[216]), .A2(n3496), .A3(MemOutputA2[248]), 
        .A4(n3317), .Y(n714) );
  OR3X1_RVT U930 ( .A1(n718), .A2(n719), .A3(n720), .Y(ipA2[23]) );
  AO221X1_RVT U931 ( .A1(MemOutputA2[23]), .A2(n3298), .A3(MemOutputA2[55]), 
        .A4(n3557), .A5(n721), .Y(n720) );
  AO22X1_RVT U932 ( .A1(MemOutputA2[87]), .A2(n3536), .A3(MemOutputA2[119]), 
        .A4(n3510), .Y(n721) );
  AO22X1_RVT U933 ( .A1(MemOutputA2[183]), .A2(n3249), .A3(MemOutputA2[151]), 
        .A4(n3283), .Y(n719) );
  AO22X1_RVT U934 ( .A1(MemOutputA2[215]), .A2(n3496), .A3(MemOutputA2[247]), 
        .A4(n3310), .Y(n718) );
  OR3X1_RVT U935 ( .A1(n722), .A2(n723), .A3(n724), .Y(ipA2[22]) );
  AO221X1_RVT U936 ( .A1(MemOutputA2[22]), .A2(n3297), .A3(MemOutputA2[54]), 
        .A4(n3557), .A5(n725), .Y(n724) );
  AO22X1_RVT U937 ( .A1(MemOutputA2[86]), .A2(n3536), .A3(MemOutputA2[118]), 
        .A4(n3509), .Y(n725) );
  AO22X1_RVT U938 ( .A1(MemOutputA2[182]), .A2(n3259), .A3(MemOutputA2[150]), 
        .A4(n3283), .Y(n723) );
  AO22X1_RVT U939 ( .A1(MemOutputA2[214]), .A2(n3496), .A3(MemOutputA2[246]), 
        .A4(n3313), .Y(n722) );
  OR3X1_RVT U940 ( .A1(n726), .A2(n727), .A3(n728), .Y(ipA2[21]) );
  AO221X1_RVT U941 ( .A1(MemOutputA2[21]), .A2(n3297), .A3(MemOutputA2[53]), 
        .A4(n3557), .A5(n729), .Y(n728) );
  AO22X1_RVT U942 ( .A1(MemOutputA2[85]), .A2(n3536), .A3(MemOutputA2[117]), 
        .A4(n3518), .Y(n729) );
  AO22X1_RVT U943 ( .A1(MemOutputA2[181]), .A2(n3254), .A3(MemOutputA2[149]), 
        .A4(n3286), .Y(n727) );
  AO22X1_RVT U944 ( .A1(MemOutputA2[213]), .A2(n3496), .A3(MemOutputA2[245]), 
        .A4(n3320), .Y(n726) );
  OR3X1_RVT U945 ( .A1(n730), .A2(n731), .A3(n732), .Y(ipA2[20]) );
  AO221X1_RVT U946 ( .A1(MemOutputA2[20]), .A2(n3298), .A3(MemOutputA2[52]), 
        .A4(n3557), .A5(n733), .Y(n732) );
  AO22X1_RVT U947 ( .A1(MemOutputA2[84]), .A2(n3536), .A3(MemOutputA2[116]), 
        .A4(n3512), .Y(n733) );
  AO22X1_RVT U949 ( .A1(MemOutputA2[212]), .A2(n3496), .A3(MemOutputA2[244]), 
        .A4(n3312), .Y(n730) );
  OR3X1_RVT U950 ( .A1(n734), .A2(n735), .A3(n736), .Y(ipA2[1]) );
  AO221X1_RVT U951 ( .A1(MemOutputA2[1]), .A2(n3307), .A3(MemOutputA2[33]), 
        .A4(n3558), .A5(n737), .Y(n736) );
  AO22X1_RVT U952 ( .A1(MemOutputA2[65]), .A2(n3537), .A3(MemOutputA2[97]), 
        .A4(n3519), .Y(n737) );
  AO22X1_RVT U953 ( .A1(MemOutputA2[161]), .A2(n3260), .A3(MemOutputA2[129]), 
        .A4(n506), .Y(n735) );
  AO22X1_RVT U954 ( .A1(MemOutputA2[193]), .A2(n3497), .A3(MemOutputA2[225]), 
        .A4(n3329), .Y(n734) );
  OR3X1_RVT U955 ( .A1(n738), .A2(n739), .A3(n740), .Y(ipA2[19]) );
  AO221X1_RVT U956 ( .A1(MemOutputA2[19]), .A2(n3297), .A3(MemOutputA2[51]), 
        .A4(n3558), .A5(n741), .Y(n740) );
  AO22X1_RVT U957 ( .A1(MemOutputA2[83]), .A2(n3537), .A3(MemOutputA2[115]), 
        .A4(n3519), .Y(n741) );
  AO22X1_RVT U958 ( .A1(MemOutputA2[179]), .A2(n3259), .A3(MemOutputA2[147]), 
        .A4(n3273), .Y(n739) );
  AO22X1_RVT U959 ( .A1(MemOutputA2[211]), .A2(n3497), .A3(MemOutputA2[243]), 
        .A4(n3326), .Y(n738) );
  OR3X1_RVT U960 ( .A1(n742), .A2(n743), .A3(n744), .Y(ipA2[18]) );
  AO221X1_RVT U961 ( .A1(MemOutputA2[18]), .A2(n3305), .A3(MemOutputA2[50]), 
        .A4(n3558), .A5(n745), .Y(n744) );
  AO22X1_RVT U962 ( .A1(MemOutputA2[82]), .A2(n3537), .A3(MemOutputA2[114]), 
        .A4(n3519), .Y(n745) );
  AO22X1_RVT U963 ( .A1(MemOutputA2[178]), .A2(n3252), .A3(MemOutputA2[146]), 
        .A4(n454), .Y(n743) );
  AO22X1_RVT U964 ( .A1(MemOutputA2[210]), .A2(n3497), .A3(MemOutputA2[242]), 
        .A4(n3325), .Y(n742) );
  OR3X1_RVT U965 ( .A1(n746), .A2(n747), .A3(n748), .Y(ipA2[17]) );
  AO221X1_RVT U966 ( .A1(MemOutputA2[17]), .A2(n3297), .A3(MemOutputA2[49]), 
        .A4(n3558), .A5(n749), .Y(n748) );
  AO22X1_RVT U967 ( .A1(MemOutputA2[81]), .A2(n3537), .A3(MemOutputA2[113]), 
        .A4(n3519), .Y(n749) );
  AO22X1_RVT U968 ( .A1(MemOutputA2[177]), .A2(n3264), .A3(MemOutputA2[145]), 
        .A4(n506), .Y(n747) );
  AO22X1_RVT U969 ( .A1(MemOutputA2[209]), .A2(n3497), .A3(MemOutputA2[241]), 
        .A4(n3330), .Y(n746) );
  OR3X1_RVT U970 ( .A1(n750), .A2(n751), .A3(n752), .Y(ipA2[16]) );
  AO221X1_RVT U971 ( .A1(MemOutputA2[16]), .A2(n3297), .A3(MemOutputA2[48]), 
        .A4(n3558), .A5(n753), .Y(n752) );
  AO22X1_RVT U972 ( .A1(MemOutputA2[80]), .A2(n3537), .A3(MemOutputA2[112]), 
        .A4(n3519), .Y(n753) );
  AO22X1_RVT U973 ( .A1(MemOutputA2[176]), .A2(n3262), .A3(MemOutputA2[144]), 
        .A4(n452), .Y(n751) );
  AO22X1_RVT U974 ( .A1(MemOutputA2[208]), .A2(n3497), .A3(MemOutputA2[240]), 
        .A4(n3322), .Y(n750) );
  OR3X1_RVT U975 ( .A1(n754), .A2(n755), .A3(n756), .Y(ipA2[15]) );
  AO221X1_RVT U976 ( .A1(MemOutputA2[15]), .A2(n3297), .A3(MemOutputA2[47]), 
        .A4(n3558), .A5(n757), .Y(n756) );
  AO22X1_RVT U977 ( .A1(MemOutputA2[79]), .A2(n3537), .A3(MemOutputA2[111]), 
        .A4(n3519), .Y(n757) );
  AO22X1_RVT U978 ( .A1(MemOutputA2[175]), .A2(n3256), .A3(MemOutputA2[143]), 
        .A4(n3282), .Y(n755) );
  AO22X1_RVT U979 ( .A1(MemOutputA2[207]), .A2(n3497), .A3(MemOutputA2[239]), 
        .A4(n3323), .Y(n754) );
  OR3X1_RVT U980 ( .A1(n758), .A2(n759), .A3(n760), .Y(ipA2[14]) );
  AO221X1_RVT U981 ( .A1(MemOutputA2[14]), .A2(n3303), .A3(MemOutputA2[46]), 
        .A4(n3558), .A5(n761), .Y(n760) );
  AO22X1_RVT U982 ( .A1(MemOutputA2[78]), .A2(n3537), .A3(MemOutputA2[110]), 
        .A4(n3519), .Y(n761) );
  AO22X1_RVT U983 ( .A1(MemOutputA2[174]), .A2(n514), .A3(MemOutputA2[142]), 
        .A4(n3285), .Y(n759) );
  AO22X1_RVT U984 ( .A1(MemOutputA2[206]), .A2(n3497), .A3(MemOutputA2[238]), 
        .A4(n3326), .Y(n758) );
  OR3X1_RVT U985 ( .A1(n762), .A2(n763), .A3(n764), .Y(ipA2[13]) );
  AO221X1_RVT U986 ( .A1(MemOutputA2[13]), .A2(n3296), .A3(MemOutputA2[45]), 
        .A4(n3558), .A5(n765), .Y(n764) );
  AO22X1_RVT U987 ( .A1(MemOutputA2[77]), .A2(n3537), .A3(MemOutputA2[109]), 
        .A4(n3519), .Y(n765) );
  AO22X1_RVT U988 ( .A1(MemOutputA2[173]), .A2(n3262), .A3(MemOutputA2[141]), 
        .A4(n454), .Y(n763) );
  AO22X1_RVT U989 ( .A1(MemOutputA2[205]), .A2(n3497), .A3(MemOutputA2[237]), 
        .A4(n3322), .Y(n762) );
  OR3X1_RVT U990 ( .A1(n766), .A2(n767), .A3(n768), .Y(ipA2[12]) );
  AO221X1_RVT U991 ( .A1(MemOutputA2[12]), .A2(n3295), .A3(MemOutputA2[44]), 
        .A4(n3558), .A5(n769), .Y(n768) );
  AO22X1_RVT U992 ( .A1(MemOutputA2[76]), .A2(n3537), .A3(MemOutputA2[108]), 
        .A4(n3519), .Y(n769) );
  AO22X1_RVT U993 ( .A1(MemOutputA2[172]), .A2(n3247), .A3(MemOutputA2[140]), 
        .A4(n3285), .Y(n767) );
  AO22X1_RVT U994 ( .A1(MemOutputA2[204]), .A2(n3497), .A3(MemOutputA2[236]), 
        .A4(n3314), .Y(n766) );
  OR3X1_RVT U995 ( .A1(n770), .A2(n771), .A3(n772), .Y(ipA2[11]) );
  AO221X1_RVT U996 ( .A1(MemOutputA2[11]), .A2(n3303), .A3(MemOutputA2[43]), 
        .A4(n3558), .A5(n773), .Y(n772) );
  AO22X1_RVT U997 ( .A1(MemOutputA2[75]), .A2(n3537), .A3(MemOutputA2[107]), 
        .A4(n3519), .Y(n773) );
  AO22X1_RVT U998 ( .A1(MemOutputA2[171]), .A2(n3250), .A3(MemOutputA2[139]), 
        .A4(n3273), .Y(n771) );
  AO22X1_RVT U999 ( .A1(MemOutputA2[203]), .A2(n3497), .A3(MemOutputA2[235]), 
        .A4(n3313), .Y(n770) );
  OR3X1_RVT U1000 ( .A1(n774), .A2(n775), .A3(n776), .Y(ipA2[10]) );
  AO221X1_RVT U1001 ( .A1(MemOutputA2[10]), .A2(n3297), .A3(MemOutputA2[42]), 
        .A4(n3558), .A5(n777), .Y(n776) );
  AO22X1_RVT U1002 ( .A1(MemOutputA2[74]), .A2(n3537), .A3(MemOutputA2[106]), 
        .A4(n3519), .Y(n777) );
  AO22X1_RVT U1003 ( .A1(MemOutputA2[170]), .A2(n451), .A3(MemOutputA2[138]), 
        .A4(n3283), .Y(n775) );
  AO22X1_RVT U1004 ( .A1(MemOutputA2[202]), .A2(n3497), .A3(MemOutputA2[234]), 
        .A4(n3310), .Y(n774) );
  OR3X1_RVT U1005 ( .A1(n778), .A2(n779), .A3(n780), .Y(ipA2[0]) );
  AO221X1_RVT U1006 ( .A1(MemOutputA2[0]), .A2(n3303), .A3(MemOutputA2[32]), 
        .A4(n3558), .A5(n781), .Y(n780) );
  AO22X1_RVT U1007 ( .A1(MemOutputA2[64]), .A2(n3537), .A3(MemOutputA2[96]), 
        .A4(n3519), .Y(n781) );
  AO22X1_RVT U1008 ( .A1(MemOutputA2[160]), .A2(n3248), .A3(MemOutputA2[128]), 
        .A4(n3272), .Y(n779) );
  OR3X1_RVT U1010 ( .A1(n782), .A2(n783), .A3(n784), .Y(ipA1[9]) );
  AO221X1_RVT U1011 ( .A1(MemOutputA1[9]), .A2(n3305), .A3(MemOutputA1[41]), 
        .A4(n3559), .A5(n785), .Y(n784) );
  AO22X1_RVT U1012 ( .A1(MemOutputA1[73]), .A2(n3538), .A3(MemOutputA1[105]), 
        .A4(n3520), .Y(n785) );
  AO22X1_RVT U1014 ( .A1(MemOutputA1[201]), .A2(n3498), .A3(MemOutputA1[233]), 
        .A4(n3310), .Y(n782) );
  OR3X1_RVT U1015 ( .A1(n786), .A2(n787), .A3(n788), .Y(ipA1[8]) );
  AO221X1_RVT U1016 ( .A1(MemOutputA1[8]), .A2(n3304), .A3(MemOutputA1[40]), 
        .A4(n3559), .A5(n789), .Y(n788) );
  AO22X1_RVT U1017 ( .A1(MemOutputA1[72]), .A2(n3538), .A3(MemOutputA1[104]), 
        .A4(n3520), .Y(n789) );
  AO22X1_RVT U1018 ( .A1(MemOutputA1[168]), .A2(n3249), .A3(MemOutputA1[136]), 
        .A4(n3270), .Y(n787) );
  AO22X1_RVT U1019 ( .A1(MemOutputA1[200]), .A2(n3498), .A3(MemOutputA1[232]), 
        .A4(n3310), .Y(n786) );
  OR3X1_RVT U1020 ( .A1(n790), .A2(n791), .A3(n792), .Y(ipA1[7]) );
  AO221X1_RVT U1021 ( .A1(MemOutputA1[7]), .A2(n3304), .A3(MemOutputA1[39]), 
        .A4(n3559), .A5(n793), .Y(n792) );
  AO22X1_RVT U1022 ( .A1(MemOutputA1[71]), .A2(n3538), .A3(MemOutputA1[103]), 
        .A4(n3520), .Y(n793) );
  AO22X1_RVT U1023 ( .A1(MemOutputA1[167]), .A2(n3263), .A3(MemOutputA1[135]), 
        .A4(n454), .Y(n791) );
  AO22X1_RVT U1024 ( .A1(MemOutputA1[199]), .A2(n3498), .A3(MemOutputA1[231]), 
        .A4(n3333), .Y(n790) );
  OR3X1_RVT U1025 ( .A1(n794), .A2(n795), .A3(n796), .Y(ipA1[6]) );
  AO221X1_RVT U1026 ( .A1(MemOutputA1[6]), .A2(n3297), .A3(MemOutputA1[38]), 
        .A4(n3559), .A5(n797), .Y(n796) );
  AO22X1_RVT U1027 ( .A1(MemOutputA1[70]), .A2(n3538), .A3(MemOutputA1[102]), 
        .A4(n3520), .Y(n797) );
  AO22X1_RVT U1028 ( .A1(MemOutputA1[166]), .A2(n451), .A3(MemOutputA1[134]), 
        .A4(n506), .Y(n795) );
  AO22X1_RVT U1029 ( .A1(MemOutputA1[198]), .A2(n3498), .A3(MemOutputA1[230]), 
        .A4(n3323), .Y(n794) );
  OR3X1_RVT U1030 ( .A1(n798), .A2(n799), .A3(n800), .Y(ipA1[5]) );
  AO221X1_RVT U1031 ( .A1(MemOutputA1[5]), .A2(n3296), .A3(MemOutputA1[37]), 
        .A4(n3559), .A5(n801), .Y(n800) );
  AO22X1_RVT U1032 ( .A1(MemOutputA1[69]), .A2(n3538), .A3(MemOutputA1[101]), 
        .A4(n3520), .Y(n801) );
  AO22X1_RVT U1033 ( .A1(MemOutputA1[165]), .A2(n3258), .A3(MemOutputA1[133]), 
        .A4(n3273), .Y(n799) );
  AO22X1_RVT U1034 ( .A1(MemOutputA1[197]), .A2(n3498), .A3(MemOutputA1[229]), 
        .A4(n3312), .Y(n798) );
  OR3X1_RVT U1035 ( .A1(n802), .A2(n803), .A3(n804), .Y(ipA1[4]) );
  AO221X1_RVT U1036 ( .A1(MemOutputA1[4]), .A2(n3299), .A3(MemOutputA1[36]), 
        .A4(n3559), .A5(n805), .Y(n804) );
  AO22X1_RVT U1037 ( .A1(MemOutputA1[68]), .A2(n3538), .A3(MemOutputA1[100]), 
        .A4(n3520), .Y(n805) );
  AO22X1_RVT U1038 ( .A1(MemOutputA1[164]), .A2(n451), .A3(MemOutputA1[132]), 
        .A4(n454), .Y(n803) );
  AO22X1_RVT U1039 ( .A1(MemOutputA1[196]), .A2(n3498), .A3(MemOutputA1[228]), 
        .A4(n3330), .Y(n802) );
  OR3X1_RVT U1040 ( .A1(n806), .A2(n807), .A3(n808), .Y(ipA1[3]) );
  AO221X1_RVT U1041 ( .A1(MemOutputA1[3]), .A2(n3298), .A3(MemOutputA1[35]), 
        .A4(n3559), .A5(n809), .Y(n808) );
  AO22X1_RVT U1042 ( .A1(MemOutputA1[67]), .A2(n3538), .A3(MemOutputA1[99]), 
        .A4(n3520), .Y(n809) );
  AO22X1_RVT U1043 ( .A1(MemOutputA1[163]), .A2(n3249), .A3(MemOutputA1[131]), 
        .A4(n454), .Y(n807) );
  AO22X1_RVT U1044 ( .A1(MemOutputA1[195]), .A2(n3498), .A3(MemOutputA1[227]), 
        .A4(n3334), .Y(n806) );
  OR3X1_RVT U1045 ( .A1(n810), .A2(n811), .A3(n812), .Y(ipA1[31]) );
  AO221X1_RVT U1046 ( .A1(MemOutputA1[31]), .A2(n3299), .A3(MemOutputA1[63]), 
        .A4(n3559), .A5(n813), .Y(n812) );
  AO22X1_RVT U1047 ( .A1(MemOutputA1[95]), .A2(n3538), .A3(MemOutputA1[127]), 
        .A4(n3520), .Y(n813) );
  AO22X1_RVT U1048 ( .A1(MemOutputA1[191]), .A2(n3252), .A3(MemOutputA1[159]), 
        .A4(n3283), .Y(n811) );
  AO22X1_RVT U1049 ( .A1(MemOutputA1[223]), .A2(n3498), .A3(MemOutputA1[255]), 
        .A4(n3324), .Y(n810) );
  OR3X1_RVT U1050 ( .A1(n814), .A2(n815), .A3(n816), .Y(ipA1[30]) );
  AO221X1_RVT U1051 ( .A1(MemOutputA1[30]), .A2(n3298), .A3(MemOutputA1[62]), 
        .A4(n3559), .A5(n817), .Y(n816) );
  AO22X1_RVT U1052 ( .A1(MemOutputA1[94]), .A2(n3538), .A3(MemOutputA1[126]), 
        .A4(n3520), .Y(n817) );
  AO22X1_RVT U1053 ( .A1(MemOutputA1[190]), .A2(n3248), .A3(MemOutputA1[158]), 
        .A4(n3276), .Y(n815) );
  AO22X1_RVT U1054 ( .A1(MemOutputA1[222]), .A2(n3498), .A3(MemOutputA1[254]), 
        .A4(n3332), .Y(n814) );
  OR3X1_RVT U1055 ( .A1(n818), .A2(n819), .A3(n820), .Y(ipA1[2]) );
  AO221X1_RVT U1056 ( .A1(MemOutputA1[2]), .A2(n3298), .A3(MemOutputA1[34]), 
        .A4(n3559), .A5(n821), .Y(n820) );
  AO22X1_RVT U1057 ( .A1(MemOutputA1[66]), .A2(n3538), .A3(MemOutputA1[98]), 
        .A4(n3520), .Y(n821) );
  AO22X1_RVT U1058 ( .A1(MemOutputA1[162]), .A2(n514), .A3(MemOutputA1[130]), 
        .A4(n3276), .Y(n819) );
  AO22X1_RVT U1059 ( .A1(MemOutputA1[194]), .A2(n3498), .A3(MemOutputA1[226]), 
        .A4(n3330), .Y(n818) );
  OR3X1_RVT U1060 ( .A1(n822), .A2(n823), .A3(n824), .Y(ipA1[29]) );
  AO221X1_RVT U1061 ( .A1(MemOutputA1[29]), .A2(n3297), .A3(MemOutputA1[61]), 
        .A4(n3559), .A5(n825), .Y(n824) );
  AO22X1_RVT U1062 ( .A1(MemOutputA1[93]), .A2(n3538), .A3(MemOutputA1[125]), 
        .A4(n3520), .Y(n825) );
  AO22X1_RVT U1063 ( .A1(MemOutputA1[189]), .A2(n514), .A3(MemOutputA1[157]), 
        .A4(n454), .Y(n823) );
  AO22X1_RVT U1064 ( .A1(MemOutputA1[221]), .A2(n3498), .A3(MemOutputA1[253]), 
        .A4(n3329), .Y(n822) );
  OR3X1_RVT U1065 ( .A1(n826), .A2(n827), .A3(n828), .Y(ipA1[28]) );
  AO221X1_RVT U1066 ( .A1(MemOutputA1[28]), .A2(n3304), .A3(MemOutputA1[60]), 
        .A4(n3559), .A5(n829), .Y(n828) );
  AO22X1_RVT U1067 ( .A1(MemOutputA1[92]), .A2(n3538), .A3(MemOutputA1[124]), 
        .A4(n3520), .Y(n829) );
  AO22X1_RVT U1068 ( .A1(MemOutputA1[188]), .A2(n3248), .A3(MemOutputA1[156]), 
        .A4(n3272), .Y(n827) );
  AO22X1_RVT U1069 ( .A1(MemOutputA1[220]), .A2(n3498), .A3(MemOutputA1[252]), 
        .A4(n3325), .Y(n826) );
  OR3X1_RVT U1070 ( .A1(n830), .A2(n831), .A3(n832), .Y(ipA1[27]) );
  AO221X1_RVT U1071 ( .A1(MemOutputA1[27]), .A2(n3297), .A3(MemOutputA1[59]), 
        .A4(n3560), .A5(n833), .Y(n832) );
  AO22X1_RVT U1072 ( .A1(MemOutputA1[91]), .A2(n519), .A3(MemOutputA1[123]), 
        .A4(n3289), .Y(n833) );
  AO22X1_RVT U1074 ( .A1(MemOutputA1[219]), .A2(n3499), .A3(MemOutputA1[251]), 
        .A4(n3312), .Y(n830) );
  OR3X1_RVT U1075 ( .A1(n834), .A2(n835), .A3(n836), .Y(ipA1[26]) );
  AO221X1_RVT U1076 ( .A1(MemOutputA1[26]), .A2(n3303), .A3(MemOutputA1[58]), 
        .A4(n3560), .A5(n837), .Y(n836) );
  AO22X1_RVT U1077 ( .A1(MemOutputA1[90]), .A2(n507), .A3(MemOutputA1[122]), 
        .A4(n3521), .Y(n837) );
  AO22X1_RVT U1078 ( .A1(MemOutputA1[186]), .A2(n3264), .A3(MemOutputA1[154]), 
        .A4(n3278), .Y(n835) );
  AO22X1_RVT U1079 ( .A1(MemOutputA1[218]), .A2(n3499), .A3(MemOutputA1[250]), 
        .A4(n3313), .Y(n834) );
  OR3X1_RVT U1080 ( .A1(n838), .A2(n839), .A3(n840), .Y(ipA1[25]) );
  AO221X1_RVT U1081 ( .A1(MemOutputA1[25]), .A2(n3307), .A3(MemOutputA1[57]), 
        .A4(n3560), .A5(n841), .Y(n840) );
  AO22X1_RVT U1082 ( .A1(MemOutputA1[89]), .A2(n519), .A3(MemOutputA1[121]), 
        .A4(n3510), .Y(n841) );
  AO22X1_RVT U1083 ( .A1(MemOutputA1[185]), .A2(n3249), .A3(MemOutputA1[153]), 
        .A4(n454), .Y(n839) );
  AO22X1_RVT U1084 ( .A1(MemOutputA1[217]), .A2(n3499), .A3(MemOutputA1[249]), 
        .A4(n3334), .Y(n838) );
  OR3X1_RVT U1085 ( .A1(n842), .A2(n843), .A3(n844), .Y(ipA1[24]) );
  AO221X1_RVT U1086 ( .A1(MemOutputA1[24]), .A2(n3307), .A3(MemOutputA1[56]), 
        .A4(n3560), .A5(n845), .Y(n844) );
  AO22X1_RVT U1087 ( .A1(MemOutputA1[88]), .A2(n507), .A3(MemOutputA1[120]), 
        .A4(n3289), .Y(n845) );
  AO22X1_RVT U1088 ( .A1(MemOutputA1[184]), .A2(n3252), .A3(MemOutputA1[152]), 
        .A4(n3283), .Y(n843) );
  AO22X1_RVT U1089 ( .A1(MemOutputA1[216]), .A2(n3499), .A3(MemOutputA1[248]), 
        .A4(n3324), .Y(n842) );
  OR3X1_RVT U1090 ( .A1(n846), .A2(n847), .A3(n848), .Y(ipA1[23]) );
  AO221X1_RVT U1091 ( .A1(MemOutputA1[23]), .A2(n3303), .A3(MemOutputA1[55]), 
        .A4(n3560), .A5(n849), .Y(n848) );
  AO22X1_RVT U1092 ( .A1(MemOutputA1[87]), .A2(n519), .A3(MemOutputA1[119]), 
        .A4(n3510), .Y(n849) );
  AO22X1_RVT U1093 ( .A1(MemOutputA1[183]), .A2(n3261), .A3(MemOutputA1[151]), 
        .A4(n506), .Y(n847) );
  AO22X1_RVT U1094 ( .A1(MemOutputA1[215]), .A2(n3499), .A3(MemOutputA1[247]), 
        .A4(n3332), .Y(n846) );
  OR3X1_RVT U1095 ( .A1(n850), .A2(n851), .A3(n852), .Y(ipA1[22]) );
  AO221X1_RVT U1096 ( .A1(MemOutputA1[22]), .A2(n3304), .A3(MemOutputA1[54]), 
        .A4(n3560), .A5(n853), .Y(n852) );
  AO22X1_RVT U1097 ( .A1(MemOutputA1[86]), .A2(n3541), .A3(MemOutputA1[118]), 
        .A4(n3289), .Y(n853) );
  AO22X1_RVT U1098 ( .A1(MemOutputA1[182]), .A2(n3260), .A3(MemOutputA1[150]), 
        .A4(n3272), .Y(n851) );
  AO22X1_RVT U1099 ( .A1(MemOutputA1[214]), .A2(n3499), .A3(MemOutputA1[246]), 
        .A4(n3332), .Y(n850) );
  OR3X1_RVT U1100 ( .A1(n854), .A2(n855), .A3(n856), .Y(ipA1[21]) );
  AO221X1_RVT U1101 ( .A1(MemOutputA1[21]), .A2(n3308), .A3(MemOutputA1[53]), 
        .A4(n3560), .A5(n857), .Y(n856) );
  AO22X1_RVT U1102 ( .A1(MemOutputA1[85]), .A2(n507), .A3(MemOutputA1[117]), 
        .A4(n3510), .Y(n857) );
  AO22X1_RVT U1103 ( .A1(MemOutputA1[181]), .A2(n3259), .A3(MemOutputA1[149]), 
        .A4(n454), .Y(n855) );
  AO22X1_RVT U1104 ( .A1(MemOutputA1[213]), .A2(n3499), .A3(MemOutputA1[245]), 
        .A4(n3325), .Y(n854) );
  OR3X1_RVT U1105 ( .A1(n858), .A2(n859), .A3(n860), .Y(ipA1[20]) );
  AO221X1_RVT U1106 ( .A1(MemOutputA1[20]), .A2(n3303), .A3(MemOutputA1[52]), 
        .A4(n3560), .A5(n861), .Y(n860) );
  AO22X1_RVT U1107 ( .A1(MemOutputA1[84]), .A2(n507), .A3(MemOutputA1[116]), 
        .A4(n3289), .Y(n861) );
  AO22X1_RVT U1108 ( .A1(MemOutputA1[180]), .A2(n3265), .A3(MemOutputA1[148]), 
        .A4(n3270), .Y(n859) );
  AO22X1_RVT U1109 ( .A1(MemOutputA1[212]), .A2(n3499), .A3(MemOutputA1[244]), 
        .A4(n3333), .Y(n858) );
  OR3X1_RVT U1110 ( .A1(n862), .A2(n863), .A3(n864), .Y(ipA1[1]) );
  AO221X1_RVT U1111 ( .A1(MemOutputA1[1]), .A2(n3299), .A3(MemOutputA1[33]), 
        .A4(n3560), .A5(n865), .Y(n864) );
  AO22X1_RVT U1112 ( .A1(MemOutputA1[65]), .A2(n3541), .A3(MemOutputA1[97]), 
        .A4(n3512), .Y(n865) );
  AO22X1_RVT U1113 ( .A1(MemOutputA1[161]), .A2(n3262), .A3(MemOutputA1[129]), 
        .A4(n3272), .Y(n863) );
  AO22X1_RVT U1114 ( .A1(MemOutputA1[193]), .A2(n3499), .A3(MemOutputA1[225]), 
        .A4(n3330), .Y(n862) );
  OR3X1_RVT U1115 ( .A1(n866), .A2(n867), .A3(n868), .Y(ipA1[19]) );
  AO221X1_RVT U1116 ( .A1(MemOutputA1[19]), .A2(n3298), .A3(MemOutputA1[51]), 
        .A4(n3560), .A5(n869), .Y(n868) );
  AO22X1_RVT U1117 ( .A1(MemOutputA1[83]), .A2(n507), .A3(MemOutputA1[115]), 
        .A4(n3510), .Y(n869) );
  AO22X1_RVT U1118 ( .A1(MemOutputA1[179]), .A2(n3257), .A3(MemOutputA1[147]), 
        .A4(n3285), .Y(n867) );
  AO22X1_RVT U1119 ( .A1(MemOutputA1[211]), .A2(n3499), .A3(MemOutputA1[243]), 
        .A4(n3334), .Y(n866) );
  OR3X1_RVT U1120 ( .A1(n870), .A2(n871), .A3(n872), .Y(ipA1[18]) );
  AO221X1_RVT U1121 ( .A1(MemOutputA1[18]), .A2(n3298), .A3(MemOutputA1[50]), 
        .A4(n3560), .A5(n873), .Y(n872) );
  AO22X1_RVT U1122 ( .A1(MemOutputA1[82]), .A2(n3541), .A3(MemOutputA1[114]), 
        .A4(n3510), .Y(n873) );
  AO22X1_RVT U1123 ( .A1(MemOutputA1[178]), .A2(n3263), .A3(MemOutputA1[146]), 
        .A4(n3281), .Y(n871) );
  AO22X1_RVT U1124 ( .A1(MemOutputA1[210]), .A2(n3499), .A3(MemOutputA1[242]), 
        .A4(n3332), .Y(n870) );
  OR3X1_RVT U1125 ( .A1(n874), .A2(n875), .A3(n876), .Y(ipA1[17]) );
  AO221X1_RVT U1126 ( .A1(MemOutputA1[17]), .A2(n3297), .A3(MemOutputA1[49]), 
        .A4(n3560), .A5(n877), .Y(n876) );
  AO22X1_RVT U1127 ( .A1(MemOutputA1[81]), .A2(n3536), .A3(MemOutputA1[113]), 
        .A4(n3289), .Y(n877) );
  AO22X1_RVT U1128 ( .A1(MemOutputA1[177]), .A2(n3249), .A3(MemOutputA1[145]), 
        .A4(n454), .Y(n875) );
  AO22X1_RVT U1129 ( .A1(MemOutputA1[209]), .A2(n3499), .A3(MemOutputA1[241]), 
        .A4(n3327), .Y(n874) );
  OR3X1_RVT U1130 ( .A1(n878), .A2(n879), .A3(n880), .Y(ipA1[16]) );
  AO221X1_RVT U1131 ( .A1(MemOutputA1[16]), .A2(n3298), .A3(MemOutputA1[48]), 
        .A4(n3561), .A5(n881), .Y(n880) );
  AO22X1_RVT U1132 ( .A1(MemOutputA1[80]), .A2(n3537), .A3(MemOutputA1[112]), 
        .A4(n3510), .Y(n881) );
  AO22X1_RVT U1133 ( .A1(MemOutputA1[176]), .A2(n3249), .A3(MemOutputA1[144]), 
        .A4(n3271), .Y(n879) );
  AO22X1_RVT U1134 ( .A1(MemOutputA1[208]), .A2(n3500), .A3(MemOutputA1[240]), 
        .A4(n3316), .Y(n878) );
  OR3X1_RVT U1135 ( .A1(n882), .A2(n883), .A3(n884), .Y(ipA1[15]) );
  AO221X1_RVT U1136 ( .A1(MemOutputA1[15]), .A2(n3298), .A3(MemOutputA1[47]), 
        .A4(n3561), .A5(n885), .Y(n884) );
  AO22X1_RVT U1137 ( .A1(MemOutputA1[79]), .A2(n507), .A3(MemOutputA1[111]), 
        .A4(n3510), .Y(n885) );
  AO22X1_RVT U1138 ( .A1(MemOutputA1[175]), .A2(n3259), .A3(MemOutputA1[143]), 
        .A4(n3286), .Y(n883) );
  AO22X1_RVT U1139 ( .A1(MemOutputA1[207]), .A2(n3500), .A3(MemOutputA1[239]), 
        .A4(n3314), .Y(n882) );
  OR3X1_RVT U1140 ( .A1(n886), .A2(n887), .A3(n888), .Y(ipA1[14]) );
  AO221X1_RVT U1141 ( .A1(MemOutputA1[14]), .A2(n3295), .A3(MemOutputA1[46]), 
        .A4(n3561), .A5(n889), .Y(n888) );
  AO22X1_RVT U1142 ( .A1(MemOutputA1[78]), .A2(n3539), .A3(MemOutputA1[110]), 
        .A4(n3510), .Y(n889) );
  AO22X1_RVT U1143 ( .A1(MemOutputA1[174]), .A2(n3248), .A3(MemOutputA1[142]), 
        .A4(n3275), .Y(n887) );
  AO22X1_RVT U1144 ( .A1(MemOutputA1[206]), .A2(n3500), .A3(MemOutputA1[238]), 
        .A4(n3316), .Y(n886) );
  OR3X1_RVT U1145 ( .A1(n890), .A2(n891), .A3(n892), .Y(ipA1[13]) );
  AO221X1_RVT U1146 ( .A1(MemOutputA1[13]), .A2(n3296), .A3(MemOutputA1[45]), 
        .A4(n3561), .A5(n893), .Y(n892) );
  AO22X1_RVT U1147 ( .A1(MemOutputA1[77]), .A2(n3539), .A3(MemOutputA1[109]), 
        .A4(n3289), .Y(n893) );
  AO22X1_RVT U1148 ( .A1(MemOutputA1[173]), .A2(n3251), .A3(MemOutputA1[141]), 
        .A4(n3276), .Y(n891) );
  AO22X1_RVT U1149 ( .A1(MemOutputA1[205]), .A2(n3500), .A3(MemOutputA1[237]), 
        .A4(n3317), .Y(n890) );
  OR3X1_RVT U1150 ( .A1(n894), .A2(n895), .A3(n896), .Y(ipA1[12]) );
  AO221X1_RVT U1151 ( .A1(MemOutputA1[12]), .A2(n3302), .A3(MemOutputA1[44]), 
        .A4(n3561), .A5(n897), .Y(n896) );
  AO22X1_RVT U1152 ( .A1(MemOutputA1[76]), .A2(n3534), .A3(MemOutputA1[108]), 
        .A4(n3521), .Y(n897) );
  AO22X1_RVT U1153 ( .A1(MemOutputA1[172]), .A2(n3262), .A3(MemOutputA1[140]), 
        .A4(n454), .Y(n895) );
  AO22X1_RVT U1154 ( .A1(MemOutputA1[204]), .A2(n3500), .A3(MemOutputA1[236]), 
        .A4(n3323), .Y(n894) );
  OR3X1_RVT U1155 ( .A1(n898), .A2(n899), .A3(n900), .Y(ipA1[11]) );
  AO221X1_RVT U1156 ( .A1(MemOutputA1[11]), .A2(n3303), .A3(MemOutputA1[43]), 
        .A4(n3561), .A5(n901), .Y(n900) );
  AO22X1_RVT U1157 ( .A1(MemOutputA1[75]), .A2(n519), .A3(MemOutputA1[107]), 
        .A4(n3521), .Y(n901) );
  AO22X1_RVT U1158 ( .A1(MemOutputA1[171]), .A2(n3259), .A3(MemOutputA1[139]), 
        .A4(n506), .Y(n899) );
  AO22X1_RVT U1159 ( .A1(MemOutputA1[203]), .A2(n3500), .A3(MemOutputA1[235]), 
        .A4(n3325), .Y(n898) );
  OR3X1_RVT U1160 ( .A1(n902), .A2(n903), .A3(n904), .Y(ipA1[10]) );
  AO221X1_RVT U1161 ( .A1(MemOutputA1[10]), .A2(n3308), .A3(MemOutputA1[42]), 
        .A4(n3561), .A5(n905), .Y(n904) );
  AO22X1_RVT U1162 ( .A1(MemOutputA1[74]), .A2(n3539), .A3(MemOutputA1[106]), 
        .A4(n3510), .Y(n905) );
  AO22X1_RVT U1163 ( .A1(MemOutputA1[170]), .A2(n451), .A3(MemOutputA1[138]), 
        .A4(n506), .Y(n903) );
  AO22X1_RVT U1164 ( .A1(MemOutputA1[202]), .A2(n3500), .A3(MemOutputA1[234]), 
        .A4(n3319), .Y(n902) );
  OR3X1_RVT U1165 ( .A1(n906), .A2(n907), .A3(n908), .Y(ipA1[0]) );
  AO221X1_RVT U1166 ( .A1(MemOutputA1[0]), .A2(n3297), .A3(MemOutputA1[32]), 
        .A4(n3561), .A5(n909), .Y(n908) );
  AO22X1_RVT U1167 ( .A1(MemOutputA1[64]), .A2(n3535), .A3(MemOutputA1[96]), 
        .A4(n3508), .Y(n909) );
  AO22X1_RVT U1168 ( .A1(MemOutputA1[160]), .A2(n3261), .A3(MemOutputA1[128]), 
        .A4(n506), .Y(n907) );
  OR3X1_RVT U1170 ( .A1(n910), .A2(n911), .A3(n912), .Y(ipA0[9]) );
  AO221X1_RVT U1171 ( .A1(MemOutputA0[9]), .A2(n3307), .A3(MemOutputA0[41]), 
        .A4(n3561), .A5(n913), .Y(n912) );
  AO22X1_RVT U1172 ( .A1(MemOutputA0[73]), .A2(n15), .A3(MemOutputA0[105]), 
        .A4(n3520), .Y(n913) );
  AO22X1_RVT U1173 ( .A1(MemOutputA0[169]), .A2(n451), .A3(MemOutputA0[137]), 
        .A4(n3283), .Y(n911) );
  AO22X1_RVT U1174 ( .A1(MemOutputA0[201]), .A2(n3500), .A3(MemOutputA0[233]), 
        .A4(n3327), .Y(n910) );
  AO221X1_RVT U1176 ( .A1(MemOutputA0[8]), .A2(n3307), .A3(MemOutputA0[40]), 
        .A4(n3561), .A5(n917), .Y(n916) );
  AO22X1_RVT U1177 ( .A1(MemOutputA0[72]), .A2(n3539), .A3(MemOutputA0[104]), 
        .A4(n3289), .Y(n917) );
  AO22X1_RVT U1178 ( .A1(MemOutputA0[168]), .A2(n3261), .A3(MemOutputA0[136]), 
        .A4(n3278), .Y(n915) );
  AO22X1_RVT U1179 ( .A1(MemOutputA0[200]), .A2(n3500), .A3(MemOutputA0[232]), 
        .A4(n3329), .Y(n914) );
  AO221X1_RVT U1181 ( .A1(MemOutputA0[7]), .A2(n3305), .A3(MemOutputA0[39]), 
        .A4(n3561), .A5(n921), .Y(n920) );
  AO22X1_RVT U1182 ( .A1(MemOutputA0[71]), .A2(n3541), .A3(MemOutputA0[103]), 
        .A4(n3289), .Y(n921) );
  AO22X1_RVT U1183 ( .A1(MemOutputA0[167]), .A2(n3260), .A3(MemOutputA0[135]), 
        .A4(n3271), .Y(n919) );
  AO22X1_RVT U1184 ( .A1(MemOutputA0[199]), .A2(n3500), .A3(MemOutputA0[231]), 
        .A4(n3325), .Y(n918) );
  AO221X1_RVT U1186 ( .A1(MemOutputA0[6]), .A2(n3305), .A3(MemOutputA0[38]), 
        .A4(n3561), .A5(n925), .Y(n924) );
  AO22X1_RVT U1187 ( .A1(MemOutputA0[70]), .A2(n3539), .A3(MemOutputA0[102]), 
        .A4(n3289), .Y(n925) );
  AO22X1_RVT U1188 ( .A1(MemOutputA0[166]), .A2(n3258), .A3(MemOutputA0[134]), 
        .A4(n3271), .Y(n923) );
  AO22X1_RVT U1189 ( .A1(MemOutputA0[198]), .A2(n3500), .A3(MemOutputA0[230]), 
        .A4(n3336), .Y(n922) );
  AO22X1_RVT U1192 ( .A1(MemOutputA0[69]), .A2(n3542), .A3(MemOutputA0[101]), 
        .A4(n3521), .Y(n929) );
  AO22X1_RVT U1202 ( .A1(MemOutputA0[67]), .A2(n3533), .A3(n508), .A4(
        MemOutputA0[99]), .Y(n937) );
  OR3X1_RVT U1205 ( .A1(n938), .A2(n939), .A3(n940), .Y(ipA0[31]) );
  AO221X1_RVT U1206 ( .A1(MemOutputA0[31]), .A2(n3298), .A3(MemOutputA0[63]), 
        .A4(n3550), .A5(n941), .Y(n940) );
  AO22X1_RVT U1207 ( .A1(MemOutputA0[95]), .A2(n3534), .A3(MemOutputA0[127]), 
        .A4(n3512), .Y(n941) );
  AO22X1_RVT U1208 ( .A1(MemOutputA0[191]), .A2(n3248), .A3(MemOutputA0[159]), 
        .A4(n3271), .Y(n939) );
  AO22X1_RVT U1209 ( .A1(MemOutputA0[223]), .A2(n3501), .A3(MemOutputA0[255]), 
        .A4(n3336), .Y(n938) );
  OR3X1_RVT U1210 ( .A1(n942), .A2(n943), .A3(n944), .Y(ipA0[30]) );
  AO221X1_RVT U1211 ( .A1(MemOutputA0[30]), .A2(n3302), .A3(MemOutputA0[62]), 
        .A4(n3560), .A5(n945), .Y(n944) );
  AO22X1_RVT U1212 ( .A1(MemOutputA0[94]), .A2(n3535), .A3(MemOutputA0[126]), 
        .A4(n3289), .Y(n945) );
  AO22X1_RVT U1213 ( .A1(MemOutputA0[190]), .A2(n3263), .A3(MemOutputA0[158]), 
        .A4(n3288), .Y(n943) );
  AO22X1_RVT U1214 ( .A1(MemOutputA0[222]), .A2(n3501), .A3(MemOutputA0[254]), 
        .A4(n3323), .Y(n942) );
  AO22X1_RVT U1217 ( .A1(n3532), .A2(MemOutputA0[66]), .A3(MemOutputA0[98]), 
        .A4(n3236), .Y(n949) );
  OR3X1_RVT U1220 ( .A1(n950), .A2(n951), .A3(n952), .Y(ipA0[29]) );
  AO221X1_RVT U1221 ( .A1(MemOutputA0[29]), .A2(n3299), .A3(MemOutputA0[61]), 
        .A4(n3558), .A5(n953), .Y(n952) );
  AO22X1_RVT U1222 ( .A1(MemOutputA0[93]), .A2(n3536), .A3(MemOutputA0[125]), 
        .A4(n3521), .Y(n953) );
  AO22X1_RVT U1223 ( .A1(MemOutputA0[189]), .A2(n3264), .A3(MemOutputA0[157]), 
        .A4(n3278), .Y(n951) );
  AO22X1_RVT U1224 ( .A1(MemOutputA0[221]), .A2(n3501), .A3(MemOutputA0[253]), 
        .A4(n3319), .Y(n950) );
  OR3X1_RVT U1225 ( .A1(n954), .A2(n955), .A3(n956), .Y(ipA0[28]) );
  AO221X1_RVT U1226 ( .A1(MemOutputA0[28]), .A2(n3298), .A3(MemOutputA0[60]), 
        .A4(n3557), .A5(n957), .Y(n956) );
  AO22X1_RVT U1227 ( .A1(MemOutputA0[92]), .A2(n3539), .A3(MemOutputA0[124]), 
        .A4(n3509), .Y(n957) );
  AO22X1_RVT U1228 ( .A1(MemOutputA0[188]), .A2(n3254), .A3(MemOutputA0[156]), 
        .A4(n454), .Y(n955) );
  AO22X1_RVT U1229 ( .A1(MemOutputA0[220]), .A2(n3501), .A3(MemOutputA0[252]), 
        .A4(n3318), .Y(n954) );
  OR3X1_RVT U1230 ( .A1(n958), .A2(n959), .A3(n960), .Y(ipA0[27]) );
  AO221X1_RVT U1231 ( .A1(MemOutputA0[27]), .A2(n3299), .A3(MemOutputA0[59]), 
        .A4(n3559), .A5(n961), .Y(n960) );
  AO22X1_RVT U1232 ( .A1(MemOutputA0[91]), .A2(n3539), .A3(MemOutputA0[123]), 
        .A4(n3517), .Y(n961) );
  AO22X1_RVT U1233 ( .A1(MemOutputA0[187]), .A2(n3253), .A3(MemOutputA0[155]), 
        .A4(n506), .Y(n959) );
  AO22X1_RVT U1234 ( .A1(MemOutputA0[219]), .A2(n3501), .A3(MemOutputA0[251]), 
        .A4(n3320), .Y(n958) );
  OR3X1_RVT U1235 ( .A1(n962), .A2(n963), .A3(n964), .Y(ipA0[26]) );
  AO221X1_RVT U1236 ( .A1(MemOutputA0[26]), .A2(n3298), .A3(MemOutputA0[58]), 
        .A4(n3546), .A5(n965), .Y(n964) );
  AO22X1_RVT U1237 ( .A1(MemOutputA0[90]), .A2(n3527), .A3(MemOutputA0[122]), 
        .A4(n3521), .Y(n965) );
  AO22X1_RVT U1238 ( .A1(MemOutputA0[186]), .A2(n3258), .A3(MemOutputA0[154]), 
        .A4(n3279), .Y(n963) );
  AO22X1_RVT U1239 ( .A1(MemOutputA0[218]), .A2(n3501), .A3(MemOutputA0[250]), 
        .A4(n3319), .Y(n962) );
  OR3X1_RVT U1240 ( .A1(n966), .A2(n967), .A3(n968), .Y(ipA0[25]) );
  AO221X1_RVT U1241 ( .A1(MemOutputA0[25]), .A2(n3298), .A3(MemOutputA0[57]), 
        .A4(n3545), .A5(n969), .Y(n968) );
  AO22X1_RVT U1242 ( .A1(MemOutputA0[89]), .A2(n3537), .A3(MemOutputA0[121]), 
        .A4(n3518), .Y(n969) );
  AO22X1_RVT U1243 ( .A1(MemOutputA0[185]), .A2(n451), .A3(MemOutputA0[153]), 
        .A4(n3273), .Y(n967) );
  AO22X1_RVT U1244 ( .A1(MemOutputA0[217]), .A2(n3501), .A3(MemOutputA0[249]), 
        .A4(n3319), .Y(n966) );
  OR3X1_RVT U1245 ( .A1(n970), .A2(n971), .A3(n972), .Y(ipA0[24]) );
  AO221X1_RVT U1246 ( .A1(MemOutputA0[24]), .A2(n3297), .A3(MemOutputA0[56]), 
        .A4(n3552), .A5(n973), .Y(n972) );
  AO22X1_RVT U1247 ( .A1(MemOutputA0[88]), .A2(n3541), .A3(MemOutputA0[120]), 
        .A4(n3508), .Y(n973) );
  AO22X1_RVT U1248 ( .A1(MemOutputA0[184]), .A2(n3248), .A3(MemOutputA0[152]), 
        .A4(n3283), .Y(n971) );
  AO22X1_RVT U1249 ( .A1(MemOutputA0[216]), .A2(n3501), .A3(MemOutputA0[248]), 
        .A4(n3317), .Y(n970) );
  OR3X1_RVT U1250 ( .A1(n974), .A2(n975), .A3(n976), .Y(ipA0[23]) );
  AO221X1_RVT U1251 ( .A1(MemOutputA0[23]), .A2(n3298), .A3(MemOutputA0[55]), 
        .A4(n3550), .A5(n977), .Y(n976) );
  AO22X1_RVT U1252 ( .A1(MemOutputA0[87]), .A2(n3531), .A3(MemOutputA0[119]), 
        .A4(n3289), .Y(n977) );
  AO22X1_RVT U1253 ( .A1(MemOutputA0[183]), .A2(n3251), .A3(MemOutputA0[151]), 
        .A4(n3285), .Y(n975) );
  AO22X1_RVT U1254 ( .A1(MemOutputA0[215]), .A2(n3496), .A3(MemOutputA0[247]), 
        .A4(n3314), .Y(n974) );
  OR3X1_RVT U1255 ( .A1(n978), .A2(n979), .A3(n980), .Y(ipA0[22]) );
  AO221X1_RVT U1256 ( .A1(MemOutputA0[22]), .A2(n3297), .A3(MemOutputA0[54]), 
        .A4(n3560), .A5(n981), .Y(n980) );
  AO22X1_RVT U1257 ( .A1(MemOutputA0[86]), .A2(n3529), .A3(MemOutputA0[118]), 
        .A4(n3519), .Y(n981) );
  AO22X1_RVT U1258 ( .A1(MemOutputA0[182]), .A2(n3264), .A3(MemOutputA0[150]), 
        .A4(n3275), .Y(n979) );
  AO22X1_RVT U1259 ( .A1(MemOutputA0[214]), .A2(n3497), .A3(MemOutputA0[246]), 
        .A4(n3315), .Y(n978) );
  OR3X1_RVT U1260 ( .A1(n982), .A2(n983), .A3(n984), .Y(ipA0[21]) );
  AO221X1_RVT U1261 ( .A1(MemOutputA0[21]), .A2(n3296), .A3(MemOutputA0[53]), 
        .A4(n3560), .A5(n985), .Y(n984) );
  AO22X1_RVT U1262 ( .A1(MemOutputA0[85]), .A2(n3530), .A3(MemOutputA0[117]), 
        .A4(n3521), .Y(n985) );
  AO22X1_RVT U1263 ( .A1(MemOutputA0[181]), .A2(n3250), .A3(MemOutputA0[149]), 
        .A4(n3276), .Y(n983) );
  AO22X1_RVT U1264 ( .A1(MemOutputA0[213]), .A2(n3496), .A3(MemOutputA0[245]), 
        .A4(n3316), .Y(n982) );
  OR3X1_RVT U1265 ( .A1(n986), .A2(n987), .A3(n988), .Y(ipA0[20]) );
  AO221X1_RVT U1266 ( .A1(MemOutputA0[20]), .A2(n3296), .A3(MemOutputA0[52]), 
        .A4(n3550), .A5(n989), .Y(n988) );
  AO22X1_RVT U1267 ( .A1(MemOutputA0[84]), .A2(n3526), .A3(MemOutputA0[116]), 
        .A4(n3506), .Y(n989) );
  AO22X1_RVT U1268 ( .A1(MemOutputA0[180]), .A2(n514), .A3(MemOutputA0[148]), 
        .A4(n3282), .Y(n987) );
  AO22X1_RVT U1269 ( .A1(MemOutputA0[212]), .A2(n3496), .A3(MemOutputA0[244]), 
        .A4(n3317), .Y(n986) );
  OR3X1_RVT U1275 ( .A1(n994), .A2(n995), .A3(n996), .Y(ipA0[19]) );
  AO221X1_RVT U1276 ( .A1(MemOutputA0[19]), .A2(n3295), .A3(MemOutputA0[51]), 
        .A4(n3550), .A5(n997), .Y(n996) );
  AO22X1_RVT U1277 ( .A1(MemOutputA0[83]), .A2(n3525), .A3(MemOutputA0[115]), 
        .A4(n3507), .Y(n997) );
  AO22X1_RVT U1278 ( .A1(MemOutputA0[179]), .A2(n3247), .A3(MemOutputA0[147]), 
        .A4(n3270), .Y(n995) );
  AO22X1_RVT U1279 ( .A1(MemOutputA0[211]), .A2(n3497), .A3(MemOutputA0[243]), 
        .A4(n3312), .Y(n994) );
  OR3X1_RVT U1280 ( .A1(n998), .A2(n999), .A3(n1000), .Y(ipA0[18]) );
  AO221X1_RVT U1281 ( .A1(MemOutputA0[18]), .A2(n3297), .A3(MemOutputA0[50]), 
        .A4(n3550), .A5(n1001), .Y(n1000) );
  AO22X1_RVT U1282 ( .A1(MemOutputA0[82]), .A2(n3543), .A3(MemOutputA0[114]), 
        .A4(n3289), .Y(n1001) );
  AO22X1_RVT U1283 ( .A1(MemOutputA0[178]), .A2(n3249), .A3(MemOutputA0[146]), 
        .A4(n3288), .Y(n999) );
  AO22X1_RVT U1284 ( .A1(MemOutputA0[210]), .A2(n3497), .A3(MemOutputA0[242]), 
        .A4(n3310), .Y(n998) );
  OR3X1_RVT U1285 ( .A1(n1002), .A2(n1003), .A3(n1004), .Y(ipA0[17]) );
  AO221X1_RVT U1286 ( .A1(MemOutputA0[17]), .A2(n3299), .A3(MemOutputA0[49]), 
        .A4(n3554), .A5(n1005), .Y(n1004) );
  AO22X1_RVT U1287 ( .A1(MemOutputA0[81]), .A2(n3543), .A3(MemOutputA0[113]), 
        .A4(n3520), .Y(n1005) );
  AO22X1_RVT U1288 ( .A1(MemOutputA0[177]), .A2(n3263), .A3(MemOutputA0[145]), 
        .A4(n3286), .Y(n1003) );
  AO22X1_RVT U1289 ( .A1(MemOutputA0[209]), .A2(n3497), .A3(MemOutputA0[241]), 
        .A4(n3320), .Y(n1002) );
  OR3X1_RVT U1290 ( .A1(n1006), .A2(n1007), .A3(n1008), .Y(ipA0[16]) );
  AO221X1_RVT U1291 ( .A1(MemOutputA0[16]), .A2(n3304), .A3(MemOutputA0[48]), 
        .A4(n3548), .A5(n1009), .Y(n1008) );
  AO22X1_RVT U1292 ( .A1(MemOutputA0[80]), .A2(n3543), .A3(MemOutputA0[112]), 
        .A4(n3521), .Y(n1009) );
  AO22X1_RVT U1294 ( .A1(MemOutputA0[208]), .A2(n3497), .A3(MemOutputA0[240]), 
        .A4(n3313), .Y(n1006) );
  OR3X1_RVT U1295 ( .A1(n1010), .A2(n1011), .A3(n1012), .Y(ipA0[15]) );
  AO221X1_RVT U1296 ( .A1(MemOutputA0[15]), .A2(n3296), .A3(MemOutputA0[47]), 
        .A4(n3551), .A5(n1013), .Y(n1012) );
  AO22X1_RVT U1297 ( .A1(MemOutputA0[79]), .A2(n3544), .A3(MemOutputA0[111]), 
        .A4(n3517), .Y(n1013) );
  AO22X1_RVT U1298 ( .A1(MemOutputA0[175]), .A2(n3248), .A3(MemOutputA0[143]), 
        .A4(n3283), .Y(n1011) );
  AO22X1_RVT U1299 ( .A1(MemOutputA0[207]), .A2(n3497), .A3(MemOutputA0[239]), 
        .A4(n3312), .Y(n1010) );
  AO221X1_RVT U1301 ( .A1(MemOutputA0[14]), .A2(n3304), .A3(MemOutputA0[46]), 
        .A4(n3549), .A5(n1017), .Y(n1016) );
  AO22X1_RVT U1302 ( .A1(MemOutputA0[78]), .A2(n3543), .A3(MemOutputA0[110]), 
        .A4(n3511), .Y(n1017) );
  AO22X1_RVT U1303 ( .A1(MemOutputA0[174]), .A2(n3265), .A3(MemOutputA0[142]), 
        .A4(n3283), .Y(n1015) );
  AO22X1_RVT U1304 ( .A1(MemOutputA0[206]), .A2(n3496), .A3(MemOutputA0[238]), 
        .A4(n3334), .Y(n1014) );
  AO221X1_RVT U1306 ( .A1(MemOutputA0[13]), .A2(n3296), .A3(MemOutputA0[45]), 
        .A4(n3547), .A5(n1021), .Y(n1020) );
  AO22X1_RVT U1307 ( .A1(MemOutputA0[77]), .A2(n3541), .A3(MemOutputA0[109]), 
        .A4(n3519), .Y(n1021) );
  AO22X1_RVT U1308 ( .A1(MemOutputA0[173]), .A2(n3259), .A3(MemOutputA0[141]), 
        .A4(n3283), .Y(n1019) );
  AO22X1_RVT U1309 ( .A1(MemOutputA0[205]), .A2(n3498), .A3(MemOutputA0[237]), 
        .A4(n3324), .Y(n1018) );
  AO221X1_RVT U1311 ( .A1(MemOutputA0[12]), .A2(n3304), .A3(MemOutputA0[44]), 
        .A4(n3549), .A5(n1025), .Y(n1024) );
  AO22X1_RVT U1312 ( .A1(MemOutputA0[76]), .A2(n3544), .A3(MemOutputA0[108]), 
        .A4(n3289), .Y(n1025) );
  AO22X1_RVT U1313 ( .A1(MemOutputA0[172]), .A2(n3257), .A3(MemOutputA0[140]), 
        .A4(n3283), .Y(n1023) );
  AO22X1_RVT U1314 ( .A1(MemOutputA0[204]), .A2(n3504), .A3(MemOutputA0[236]), 
        .A4(n3333), .Y(n1022) );
  OR3X1_RVT U1315 ( .A1(n1026), .A2(n1027), .A3(n1028), .Y(ipA0[11]) );
  AO221X1_RVT U1316 ( .A1(MemOutputA0[11]), .A2(n3304), .A3(MemOutputA0[43]), 
        .A4(n3564), .A5(n1029), .Y(n1028) );
  AO22X1_RVT U1317 ( .A1(MemOutputA0[75]), .A2(n3541), .A3(MemOutputA0[107]), 
        .A4(n3511), .Y(n1029) );
  AO22X1_RVT U1318 ( .A1(MemOutputA0[171]), .A2(n3262), .A3(MemOutputA0[139]), 
        .A4(n3276), .Y(n1027) );
  AO22X1_RVT U1319 ( .A1(MemOutputA0[203]), .A2(n3504), .A3(MemOutputA0[235]), 
        .A4(n3330), .Y(n1026) );
  AO221X1_RVT U1321 ( .A1(MemOutputA0[10]), .A2(n3303), .A3(MemOutputA0[42]), 
        .A4(n3545), .A5(n1033), .Y(n1032) );
  AO22X1_RVT U1323 ( .A1(MemOutputA0[170]), .A2(n3263), .A3(MemOutputA0[138]), 
        .A4(n3281), .Y(n1031) );
  AO22X1_RVT U1324 ( .A1(MemOutputA0[202]), .A2(n3502), .A3(MemOutputA0[234]), 
        .A4(n3332), .Y(n1030) );
  AO22X1_RVT U1327 ( .A1(n12), .A2(MemOutputA0[64]), .A3(n3514), .A4(
        MemOutputA0[96]), .Y(n1037) );
  AND2X1_RVT U1342 ( .A1(opC11_d3_6_), .A2(n3349), .Y(N999) );
  AND2X1_RVT U1343 ( .A1(opC11_out[31]), .A2(n3359), .Y(N960) );
  AND2X1_RVT U1344 ( .A1(opC11_out[30]), .A2(n3359), .Y(N959) );
  AND2X1_RVT U1345 ( .A1(opC11_out[29]), .A2(n3359), .Y(N958) );
  AND2X1_RVT U1346 ( .A1(opC11_out[28]), .A2(n3359), .Y(N957) );
  AND2X1_RVT U1347 ( .A1(opC11_out[27]), .A2(n3359), .Y(N956) );
  AND2X1_RVT U1348 ( .A1(opC11_out[26]), .A2(n3359), .Y(N955) );
  AND2X1_RVT U1349 ( .A1(opC11_out[25]), .A2(n3359), .Y(N954) );
  AND2X1_RVT U1350 ( .A1(opC11_out[24]), .A2(n3359), .Y(N953) );
  AND2X1_RVT U1351 ( .A1(opC11_out[23]), .A2(n3345), .Y(N952) );
  AND2X1_RVT U1352 ( .A1(opC11_out[22]), .A2(n3472), .Y(N951) );
  AND2X1_RVT U1353 ( .A1(opC11_out[21]), .A2(n3472), .Y(N950) );
  AND2X1_RVT U1354 ( .A1(opC11_out[20]), .A2(n3472), .Y(N949) );
  AND2X1_RVT U1355 ( .A1(opC11_out[19]), .A2(n3472), .Y(N948) );
  AND2X1_RVT U1356 ( .A1(opC11_out[18]), .A2(n3472), .Y(N947) );
  AND2X1_RVT U1357 ( .A1(opC11_out[17]), .A2(n3472), .Y(N946) );
  AND2X1_RVT U1358 ( .A1(opC11_out[16]), .A2(n3472), .Y(N945) );
  AND2X1_RVT U1359 ( .A1(opC11_out[15]), .A2(n3472), .Y(N944) );
  AND2X1_RVT U1360 ( .A1(opC11_out[14]), .A2(n3472), .Y(N943) );
  AND2X1_RVT U1361 ( .A1(opC11_out[13]), .A2(n3472), .Y(N942) );
  AND2X1_RVT U1362 ( .A1(opC11_out[12]), .A2(n3472), .Y(N941) );
  AND2X1_RVT U1363 ( .A1(opC11_out[11]), .A2(n3456), .Y(N940) );
  AND2X1_RVT U1364 ( .A1(opC11_out[10]), .A2(n3458), .Y(N939) );
  AND2X1_RVT U1365 ( .A1(opC11_out[9]), .A2(n3459), .Y(N938) );
  AND2X1_RVT U1366 ( .A1(opC11_out[8]), .A2(n3460), .Y(N937) );
  AND2X1_RVT U1367 ( .A1(opC11_out[7]), .A2(n3441), .Y(N936) );
  AND2X1_RVT U1368 ( .A1(opC11_out[6]), .A2(n3464), .Y(N935) );
  AND2X1_RVT U1369 ( .A1(opC11_out[5]), .A2(n3474), .Y(N934) );
  AND2X1_RVT U1370 ( .A1(opC11_out[4]), .A2(n3476), .Y(N933) );
  AND2X1_RVT U1371 ( .A1(opC11_out[3]), .A2(n3475), .Y(N932) );
  AND2X1_RVT U1372 ( .A1(opC11_out[2]), .A2(n3441), .Y(N931) );
  AND2X1_RVT U1373 ( .A1(opC11_out[1]), .A2(n3441), .Y(N930) );
  AND2X1_RVT U1375 ( .A1(opC02_out[31]), .A2(n3343), .Y(N832) );
  AND2X1_RVT U1376 ( .A1(opC02_out[30]), .A2(n3343), .Y(N831) );
  AND2X1_RVT U1377 ( .A1(opC02_out[29]), .A2(n3343), .Y(N830) );
  AND2X1_RVT U1378 ( .A1(opC02_out[28]), .A2(n3343), .Y(N829) );
  AND2X1_RVT U1379 ( .A1(opC02_out[27]), .A2(n3343), .Y(N828) );
  AND2X1_RVT U1380 ( .A1(opC02_out[26]), .A2(n3343), .Y(N827) );
  AND2X1_RVT U1381 ( .A1(opC02_out[25]), .A2(n3343), .Y(N826) );
  AND2X1_RVT U1382 ( .A1(opC02_out[24]), .A2(n3343), .Y(N825) );
  AND2X1_RVT U1383 ( .A1(opC02_out[23]), .A2(n3343), .Y(N824) );
  AND2X1_RVT U1384 ( .A1(opC02_out[22]), .A2(n3343), .Y(N823) );
  AND2X1_RVT U1385 ( .A1(opC02_out[21]), .A2(n3343), .Y(N822) );
  AND2X1_RVT U1386 ( .A1(opC02_out[20]), .A2(n3343), .Y(N821) );
  AND2X1_RVT U1387 ( .A1(opC02_out[19]), .A2(n3344), .Y(N820) );
  AND2X1_RVT U1388 ( .A1(opC02_out[18]), .A2(n3344), .Y(N819) );
  AND2X1_RVT U1389 ( .A1(opC02_out[17]), .A2(n3344), .Y(N818) );
  AND2X1_RVT U1390 ( .A1(opC02_out[16]), .A2(n3344), .Y(N817) );
  AND2X1_RVT U1391 ( .A1(opC02_out[15]), .A2(n3344), .Y(N816) );
  AND2X1_RVT U1392 ( .A1(opC02_out[14]), .A2(n3344), .Y(N815) );
  AND2X1_RVT U1393 ( .A1(opC02_out[13]), .A2(n3344), .Y(N814) );
  AND2X1_RVT U1394 ( .A1(opC02_out[12]), .A2(n3344), .Y(N813) );
  AND2X1_RVT U1395 ( .A1(opC02_out[11]), .A2(n3344), .Y(N812) );
  AND2X1_RVT U1396 ( .A1(opC02_out[10]), .A2(n3344), .Y(N811) );
  AND2X1_RVT U1397 ( .A1(opC02_out[9]), .A2(n3344), .Y(N810) );
  AND2X1_RVT U1398 ( .A1(opC02_out[8]), .A2(n3345), .Y(N809) );
  AND2X1_RVT U1399 ( .A1(opC02_out[7]), .A2(n3345), .Y(N808) );
  AND2X1_RVT U1400 ( .A1(opC02_out[6]), .A2(n3345), .Y(N807) );
  AND2X1_RVT U1401 ( .A1(opC02_out[5]), .A2(n3345), .Y(N806) );
  AND2X1_RVT U1402 ( .A1(opC02_out[4]), .A2(n3345), .Y(N805) );
  AND2X1_RVT U1403 ( .A1(opC02_out[3]), .A2(n3345), .Y(N804) );
  AND2X1_RVT U1404 ( .A1(opC02_out[2]), .A2(n3345), .Y(N803) );
  AND2X1_RVT U1405 ( .A1(opC02_out[1]), .A2(n3345), .Y(N802) );
  AND2X1_RVT U1406 ( .A1(opC02_out[0]), .A2(n3345), .Y(N801) );
  AND2X1_RVT U1407 ( .A1(opC10_out[31]), .A2(n3345), .Y(N672) );
  AND2X1_RVT U1408 ( .A1(opC10_out[30]), .A2(n3345), .Y(N671) );
  AND2X1_RVT U1409 ( .A1(opC10_out[29]), .A2(n3346), .Y(N670) );
  AND2X1_RVT U1410 ( .A1(opC10_out[28]), .A2(n3346), .Y(N669) );
  AND2X1_RVT U1411 ( .A1(opC10_out[27]), .A2(n3346), .Y(N668) );
  AND2X1_RVT U1412 ( .A1(opC10_out[26]), .A2(n3346), .Y(N667) );
  AND2X1_RVT U1413 ( .A1(opC10_out[25]), .A2(n3346), .Y(N666) );
  AND2X1_RVT U1414 ( .A1(opC10_out[24]), .A2(n3346), .Y(N665) );
  AND2X1_RVT U1415 ( .A1(opC10_out[23]), .A2(n3346), .Y(N664) );
  AND2X1_RVT U1416 ( .A1(opC10_out[22]), .A2(n3346), .Y(N663) );
  AND2X1_RVT U1417 ( .A1(opC10_out[21]), .A2(n3346), .Y(N662) );
  AND2X1_RVT U1418 ( .A1(opC10_out[20]), .A2(n3346), .Y(N661) );
  AND2X1_RVT U1419 ( .A1(opC10_out[19]), .A2(n3346), .Y(N660) );
  AND2X1_RVT U1420 ( .A1(opC10_out[18]), .A2(n3346), .Y(N659) );
  AND2X1_RVT U1421 ( .A1(opC10_out[17]), .A2(n3347), .Y(N658) );
  AND2X1_RVT U1422 ( .A1(opC10_out[16]), .A2(n3347), .Y(N657) );
  AND2X1_RVT U1423 ( .A1(opC10_out[15]), .A2(n3347), .Y(N656) );
  AND2X1_RVT U1424 ( .A1(opC10_out[14]), .A2(n3347), .Y(N655) );
  AND2X1_RVT U1425 ( .A1(opC10_out[13]), .A2(n3347), .Y(N654) );
  AND2X1_RVT U1426 ( .A1(opC10_out[12]), .A2(n3347), .Y(N653) );
  AND2X1_RVT U1427 ( .A1(opC10_out[11]), .A2(n3347), .Y(N652) );
  AND2X1_RVT U1428 ( .A1(opC10_out[10]), .A2(n3347), .Y(N651) );
  AND2X1_RVT U1429 ( .A1(opC10_out[9]), .A2(n3347), .Y(N650) );
  AND2X1_RVT U1430 ( .A1(opC10_out[8]), .A2(n3347), .Y(N649) );
  AND2X1_RVT U1431 ( .A1(opC10_out[7]), .A2(n3347), .Y(N648) );
  AND2X1_RVT U1432 ( .A1(opC10_out[6]), .A2(n3347), .Y(N647) );
  AND2X1_RVT U1433 ( .A1(opC10_out[5]), .A2(n3348), .Y(N646) );
  AND2X1_RVT U1434 ( .A1(opC10_out[4]), .A2(n3348), .Y(N645) );
  AND2X1_RVT U1435 ( .A1(opC10_out[3]), .A2(n3348), .Y(N644) );
  AND2X1_RVT U1436 ( .A1(opC10_out[2]), .A2(n3348), .Y(N643) );
  AND2X1_RVT U1437 ( .A1(opC10_out[1]), .A2(n3348), .Y(N642) );
  AND2X1_RVT U1438 ( .A1(opC10_out[0]), .A2(n3348), .Y(N641) );
  AND2X1_RVT U1439 ( .A1(opC01_out[31]), .A2(n3348), .Y(N512) );
  AND2X1_RVT U1440 ( .A1(opC01_out[30]), .A2(n3348), .Y(N511) );
  AND2X1_RVT U1441 ( .A1(opC01_out[29]), .A2(n3348), .Y(N510) );
  AND2X1_RVT U1442 ( .A1(opC01_out[28]), .A2(n3348), .Y(N509) );
  AND2X1_RVT U1443 ( .A1(opC01_out[27]), .A2(n3348), .Y(N508) );
  AND2X1_RVT U1444 ( .A1(opC01_out[26]), .A2(n3348), .Y(N507) );
  AND2X1_RVT U1445 ( .A1(opC01_out[25]), .A2(n3349), .Y(N506) );
  AND2X1_RVT U1446 ( .A1(opC01_out[24]), .A2(n3344), .Y(N505) );
  AND2X1_RVT U1447 ( .A1(opC01_out[23]), .A2(n3472), .Y(N504) );
  AND2X1_RVT U1448 ( .A1(opC01_out[22]), .A2(n3350), .Y(N503) );
  AND2X1_RVT U1449 ( .A1(opC01_out[21]), .A2(n3355), .Y(N502) );
  AND2X1_RVT U1450 ( .A1(opC01_out[20]), .A2(n3350), .Y(N501) );
  AND2X1_RVT U1451 ( .A1(opC01_out[19]), .A2(n3350), .Y(N500) );
  AND2X1_RVT U1452 ( .A1(opC01_out[18]), .A2(n3350), .Y(N499) );
  AND2X1_RVT U1453 ( .A1(opC01_out[17]), .A2(n3350), .Y(N498) );
  AND2X1_RVT U1454 ( .A1(opC01_out[16]), .A2(n3351), .Y(N497) );
  AND2X1_RVT U1455 ( .A1(opC01_out[15]), .A2(n3350), .Y(N496) );
  AND2X1_RVT U1456 ( .A1(opC01_out[14]), .A2(n3351), .Y(N495) );
  AND2X1_RVT U1457 ( .A1(opC01_out[13]), .A2(n3350), .Y(N494) );
  AND2X1_RVT U1458 ( .A1(opC01_out[12]), .A2(n3351), .Y(N493) );
  AND2X1_RVT U1459 ( .A1(opC01_out[11]), .A2(n3351), .Y(N492) );
  AND2X1_RVT U1460 ( .A1(opC01_out[10]), .A2(n3351), .Y(N491) );
  AND2X1_RVT U1461 ( .A1(opC01_out[9]), .A2(n3351), .Y(N490) );
  AND2X1_RVT U1462 ( .A1(opC01_out[8]), .A2(n3351), .Y(N489) );
  AND2X1_RVT U1463 ( .A1(opC01_out[7]), .A2(n3351), .Y(N488) );
  AND2X1_RVT U1464 ( .A1(opC01_out[6]), .A2(n3351), .Y(N487) );
  AND2X1_RVT U1465 ( .A1(opC01_out[5]), .A2(n3351), .Y(N486) );
  AND2X1_RVT U1466 ( .A1(opC01_out[4]), .A2(n3351), .Y(N485) );
  AND2X1_RVT U1467 ( .A1(opC01_out[3]), .A2(n3352), .Y(N484) );
  AND2X1_RVT U1468 ( .A1(opC01_out[2]), .A2(n3351), .Y(N483) );
  AND2X1_RVT U1469 ( .A1(opC01_out[1]), .A2(n3352), .Y(N482) );
  AND2X1_RVT U1470 ( .A1(opC01_out[0]), .A2(n3352), .Y(N481) );
  AND2X1_RVT U1471 ( .A1(opC32_out[31]), .A2(n3352), .Y(N1824) );
  AND2X1_RVT U1472 ( .A1(opC32_out[30]), .A2(n3352), .Y(N1823) );
  AND2X1_RVT U1473 ( .A1(opC32_out[29]), .A2(n3352), .Y(N1822) );
  AND2X1_RVT U1474 ( .A1(opC32_out[28]), .A2(n3352), .Y(N1821) );
  AND2X1_RVT U1475 ( .A1(opC32_out[27]), .A2(n3352), .Y(N1820) );
  AND2X1_RVT U1476 ( .A1(opC32_out[26]), .A2(n3352), .Y(N1819) );
  AND2X1_RVT U1477 ( .A1(opC32_out[25]), .A2(n3352), .Y(N1818) );
  AND2X1_RVT U1478 ( .A1(opC32_out[24]), .A2(n3352), .Y(N1817) );
  AND2X1_RVT U1479 ( .A1(opC32_out[23]), .A2(n3353), .Y(N1816) );
  AND2X1_RVT U1480 ( .A1(opC32_out[22]), .A2(n3352), .Y(N1815) );
  AND2X1_RVT U1481 ( .A1(opC32_out[21]), .A2(n3353), .Y(N1814) );
  AND2X1_RVT U1482 ( .A1(opC32_out[20]), .A2(n3353), .Y(N1813) );
  AND2X1_RVT U1483 ( .A1(opC32_out[19]), .A2(n3353), .Y(N1812) );
  AND2X1_RVT U1484 ( .A1(opC32_out[18]), .A2(n3353), .Y(N1811) );
  AND2X1_RVT U1485 ( .A1(opC32_out[17]), .A2(n3353), .Y(N1810) );
  AND2X1_RVT U1486 ( .A1(opC32_out[16]), .A2(n3353), .Y(N1809) );
  AND2X1_RVT U1487 ( .A1(opC32_out[15]), .A2(n3353), .Y(N1808) );
  AND2X1_RVT U1488 ( .A1(opC32_out[14]), .A2(n3353), .Y(N1807) );
  AND2X1_RVT U1489 ( .A1(opC32_out[13]), .A2(n3353), .Y(N1806) );
  AND2X1_RVT U1490 ( .A1(opC32_out[12]), .A2(n3353), .Y(N1805) );
  AND2X1_RVT U1491 ( .A1(opC32_out[11]), .A2(n3354), .Y(N1804) );
  AND2X1_RVT U1492 ( .A1(opC32_out[10]), .A2(n3353), .Y(N1803) );
  AND2X1_RVT U1493 ( .A1(opC32_out[9]), .A2(n3354), .Y(N1802) );
  AND2X1_RVT U1494 ( .A1(opC32_out[8]), .A2(n3354), .Y(N1801) );
  AND2X1_RVT U1495 ( .A1(opC32_out[7]), .A2(n3358), .Y(N1800) );
  AND2X1_RVT U1496 ( .A1(opC32_out[6]), .A2(n3354), .Y(N1799) );
  AND2X1_RVT U1497 ( .A1(opC32_out[5]), .A2(n3354), .Y(N1798) );
  AND2X1_RVT U1498 ( .A1(opC32_out[4]), .A2(n3354), .Y(N1797) );
  AND2X1_RVT U1499 ( .A1(opC32_out[3]), .A2(n3354), .Y(N1796) );
  AND2X1_RVT U1500 ( .A1(opC32_out[2]), .A2(n3354), .Y(N1795) );
  AND2X1_RVT U1501 ( .A1(opC32_out[1]), .A2(n3354), .Y(N1794) );
  AND2X1_RVT U1502 ( .A1(opC32_out[0]), .A2(n3354), .Y(N1793) );
  AND2X1_RVT U1503 ( .A1(opC23_out[31]), .A2(n3354), .Y(N1792) );
  AND2X1_RVT U1504 ( .A1(opC23_out[30]), .A2(n3355), .Y(N1791) );
  AND2X1_RVT U1505 ( .A1(opC23_out[29]), .A2(n3355), .Y(N1790) );
  AND2X1_RVT U1506 ( .A1(opC23_out[28]), .A2(n3355), .Y(N1789) );
  AND2X1_RVT U1507 ( .A1(opC23_out[27]), .A2(n3355), .Y(N1788) );
  AND2X1_RVT U1508 ( .A1(opC23_out[26]), .A2(n3355), .Y(N1787) );
  AND2X1_RVT U1509 ( .A1(opC23_out[25]), .A2(n3355), .Y(N1786) );
  AND2X1_RVT U1510 ( .A1(opC23_out[24]), .A2(n3355), .Y(N1785) );
  AND2X1_RVT U1511 ( .A1(opC23_out[23]), .A2(n3355), .Y(N1784) );
  AND2X1_RVT U1512 ( .A1(opC23_out[22]), .A2(n3355), .Y(N1783) );
  AND2X1_RVT U1513 ( .A1(opC23_out[21]), .A2(n3355), .Y(N1782) );
  AND2X1_RVT U1514 ( .A1(opC23_out[20]), .A2(n3355), .Y(N1781) );
  AND2X1_RVT U1515 ( .A1(opC23_out[19]), .A2(n3356), .Y(N1780) );
  AND2X1_RVT U1516 ( .A1(opC23_out[18]), .A2(n3356), .Y(N1779) );
  AND2X1_RVT U1517 ( .A1(opC23_out[17]), .A2(n3356), .Y(N1778) );
  AND2X1_RVT U1518 ( .A1(opC23_out[16]), .A2(n3356), .Y(N1777) );
  AND2X1_RVT U1519 ( .A1(opC23_out[15]), .A2(n3356), .Y(N1776) );
  AND2X1_RVT U1520 ( .A1(opC23_out[14]), .A2(n3356), .Y(N1775) );
  AND2X1_RVT U1521 ( .A1(opC23_out[13]), .A2(n3356), .Y(N1774) );
  AND2X1_RVT U1522 ( .A1(opC23_out[12]), .A2(n3356), .Y(N1773) );
  AND2X1_RVT U1523 ( .A1(opC23_out[11]), .A2(n3356), .Y(N1772) );
  AND2X1_RVT U1524 ( .A1(opC23_out[10]), .A2(n3356), .Y(N1771) );
  AND2X1_RVT U1525 ( .A1(opC23_out[9]), .A2(n3356), .Y(N1770) );
  AND2X1_RVT U1526 ( .A1(opC23_out[8]), .A2(n3356), .Y(N1769) );
  AND2X1_RVT U1527 ( .A1(opC23_out[7]), .A2(n3357), .Y(N1768) );
  AND2X1_RVT U1528 ( .A1(opC23_out[6]), .A2(n3357), .Y(N1767) );
  AND2X1_RVT U1529 ( .A1(opC23_out[5]), .A2(n3357), .Y(N1766) );
  AND2X1_RVT U1530 ( .A1(opC23_out[4]), .A2(n3357), .Y(N1765) );
  AND2X1_RVT U1531 ( .A1(opC23_out[3]), .A2(n3357), .Y(N1764) );
  AND2X1_RVT U1532 ( .A1(opC23_out[2]), .A2(n3357), .Y(N1763) );
  AND2X1_RVT U1533 ( .A1(opC23_out[1]), .A2(n3357), .Y(N1762) );
  AND2X1_RVT U1534 ( .A1(opC23_out[0]), .A2(n3357), .Y(N1761) );
  AND2X1_RVT U1535 ( .A1(opC31_out[31]), .A2(n3357), .Y(N1728) );
  AND2X1_RVT U1536 ( .A1(opC31_out[30]), .A2(n3354), .Y(N1727) );
  AND2X1_RVT U1537 ( .A1(opC31_out[29]), .A2(n3357), .Y(N1726) );
  AND2X1_RVT U1538 ( .A1(opC31_out[28]), .A2(n3357), .Y(N1725) );
  AND2X1_RVT U1539 ( .A1(opC31_out[27]), .A2(n3357), .Y(N1724) );
  AND2X1_RVT U1540 ( .A1(opC31_out[26]), .A2(n3358), .Y(N1723) );
  AND2X1_RVT U1541 ( .A1(opC31_out[25]), .A2(n3358), .Y(N1722) );
  AND2X1_RVT U1542 ( .A1(opC31_out[24]), .A2(n3358), .Y(N1721) );
  AND2X1_RVT U1543 ( .A1(opC31_out[23]), .A2(n3358), .Y(N1720) );
  AND2X1_RVT U1544 ( .A1(opC31_out[22]), .A2(n3358), .Y(N1719) );
  AND2X1_RVT U1545 ( .A1(opC31_out[21]), .A2(n3358), .Y(N1718) );
  AND2X1_RVT U1546 ( .A1(opC31_out[20]), .A2(n3358), .Y(N1717) );
  AND2X1_RVT U1547 ( .A1(opC31_out[19]), .A2(n3358), .Y(N1716) );
  AND2X1_RVT U1548 ( .A1(opC31_out[18]), .A2(n3358), .Y(N1715) );
  AND2X1_RVT U1549 ( .A1(opC31_out[17]), .A2(n3358), .Y(N1714) );
  AND2X1_RVT U1550 ( .A1(opC31_out[16]), .A2(n3358), .Y(N1713) );
  AND2X1_RVT U1551 ( .A1(opC31_out[15]), .A2(n3472), .Y(N1712) );
  AND2X1_RVT U1552 ( .A1(opC31_out[14]), .A2(n3464), .Y(N1711) );
  AND2X1_RVT U1553 ( .A1(opC31_out[13]), .A2(n3470), .Y(N1710) );
  AND2X1_RVT U1554 ( .A1(opC31_out[12]), .A2(n3469), .Y(N1709) );
  AND2X1_RVT U1555 ( .A1(opC31_out[11]), .A2(n3471), .Y(N1708) );
  AND2X1_RVT U1556 ( .A1(opC31_out[10]), .A2(n3468), .Y(N1707) );
  AND2X1_RVT U1557 ( .A1(opC31_out[9]), .A2(n3467), .Y(N1706) );
  AND2X1_RVT U1558 ( .A1(opC31_out[8]), .A2(n3475), .Y(N1705) );
  AND2X1_RVT U1559 ( .A1(opC31_out[7]), .A2(n3364), .Y(N1704) );
  AND2X1_RVT U1560 ( .A1(opC31_out[6]), .A2(n3359), .Y(N1703) );
  AND2X1_RVT U1561 ( .A1(opC31_out[5]), .A2(n3359), .Y(N1702) );
  AND2X1_RVT U1562 ( .A1(opC31_out[4]), .A2(n3359), .Y(N1701) );
  AND2X1_RVT U1563 ( .A1(opC31_out[3]), .A2(n3360), .Y(N1700) );
  AND2X1_RVT U1564 ( .A1(opC31_out[2]), .A2(n3360), .Y(N1699) );
  AND2X1_RVT U1565 ( .A1(opC31_out[1]), .A2(n3360), .Y(N1698) );
  AND2X1_RVT U1566 ( .A1(opC31_out[0]), .A2(n3360), .Y(N1697) );
  AND2X1_RVT U1567 ( .A1(opC22_out[31]), .A2(n3360), .Y(N1664) );
  AND2X1_RVT U1568 ( .A1(opC22_out[30]), .A2(n3360), .Y(N1663) );
  AND2X1_RVT U1569 ( .A1(opC22_out[29]), .A2(n3360), .Y(N1662) );
  AND2X1_RVT U1570 ( .A1(opC22_out[28]), .A2(n3360), .Y(N1661) );
  AND2X1_RVT U1571 ( .A1(opC22_out[27]), .A2(n3360), .Y(N1660) );
  AND2X1_RVT U1572 ( .A1(opC22_out[26]), .A2(n3360), .Y(N1659) );
  AND2X1_RVT U1573 ( .A1(opC22_out[25]), .A2(n3360), .Y(N1658) );
  AND2X1_RVT U1574 ( .A1(opC22_out[24]), .A2(n3360), .Y(N1657) );
  AND2X1_RVT U1575 ( .A1(opC22_out[23]), .A2(n3361), .Y(N1656) );
  AND2X1_RVT U1576 ( .A1(opC22_out[22]), .A2(n3361), .Y(N1655) );
  AND2X1_RVT U1577 ( .A1(opC22_out[21]), .A2(n3361), .Y(N1654) );
  AND2X1_RVT U1578 ( .A1(opC22_out[20]), .A2(n3361), .Y(N1653) );
  AND2X1_RVT U1579 ( .A1(opC22_out[19]), .A2(n3361), .Y(N1652) );
  AND2X1_RVT U1580 ( .A1(opC22_out[18]), .A2(n3361), .Y(N1651) );
  AND2X1_RVT U1581 ( .A1(opC22_out[17]), .A2(n3361), .Y(N1650) );
  AND2X1_RVT U1582 ( .A1(opC22_out[16]), .A2(n3361), .Y(N1649) );
  AND2X1_RVT U1583 ( .A1(opC22_out[15]), .A2(n3361), .Y(N1648) );
  AND2X1_RVT U1584 ( .A1(opC22_out[14]), .A2(n3361), .Y(N1647) );
  AND2X1_RVT U1585 ( .A1(opC22_out[13]), .A2(n3361), .Y(N1646) );
  AND2X1_RVT U1586 ( .A1(opC22_out[12]), .A2(n3361), .Y(N1645) );
  AND2X1_RVT U1587 ( .A1(opC22_out[11]), .A2(n3362), .Y(N1644) );
  AND2X1_RVT U1588 ( .A1(opC22_out[10]), .A2(n3362), .Y(N1643) );
  AND2X1_RVT U1589 ( .A1(opC22_out[9]), .A2(n3362), .Y(N1642) );
  AND2X1_RVT U1590 ( .A1(opC22_out[8]), .A2(n3362), .Y(N1641) );
  AND2X1_RVT U1591 ( .A1(opC22_out[7]), .A2(n3362), .Y(N1640) );
  AND2X1_RVT U1592 ( .A1(opC22_out[6]), .A2(n3362), .Y(N1639) );
  AND2X1_RVT U1593 ( .A1(opC22_out[5]), .A2(n3362), .Y(N1638) );
  AND2X1_RVT U1594 ( .A1(opC22_out[4]), .A2(n3362), .Y(N1637) );
  AND2X1_RVT U1595 ( .A1(opC22_out[3]), .A2(n3362), .Y(N1636) );
  AND2X1_RVT U1596 ( .A1(opC22_out[2]), .A2(n3362), .Y(N1635) );
  AND2X1_RVT U1597 ( .A1(opC22_out[1]), .A2(n3362), .Y(N1634) );
  AND2X1_RVT U1598 ( .A1(opC22_out[0]), .A2(n3362), .Y(N1633) );
  AND2X1_RVT U1599 ( .A1(opC13_out[31]), .A2(n3363), .Y(N1600) );
  AND2X1_RVT U1600 ( .A1(opC13_out[30]), .A2(n3363), .Y(N1599) );
  AND2X1_RVT U1601 ( .A1(opC13_out[29]), .A2(n3363), .Y(N1598) );
  AND2X1_RVT U1602 ( .A1(opC13_out[28]), .A2(n3363), .Y(N1597) );
  AND2X1_RVT U1603 ( .A1(opC13_out[27]), .A2(n3363), .Y(N1596) );
  AND2X1_RVT U1604 ( .A1(opC13_out[26]), .A2(n3363), .Y(N1595) );
  AND2X1_RVT U1605 ( .A1(opC13_out[25]), .A2(n3363), .Y(N1594) );
  AND2X1_RVT U1606 ( .A1(opC13_out[24]), .A2(n3363), .Y(N1593) );
  AND2X1_RVT U1607 ( .A1(opC13_out[23]), .A2(n3363), .Y(N1592) );
  AND2X1_RVT U1608 ( .A1(opC13_out[22]), .A2(n3363), .Y(N1591) );
  AND2X1_RVT U1609 ( .A1(opC13_out[21]), .A2(n3363), .Y(N1590) );
  AND2X1_RVT U1610 ( .A1(opC13_out[20]), .A2(n3363), .Y(N1589) );
  AND2X1_RVT U1611 ( .A1(opC13_out[19]), .A2(n3364), .Y(N1588) );
  AND2X1_RVT U1612 ( .A1(opC13_out[18]), .A2(n3364), .Y(N1587) );
  AND2X1_RVT U1613 ( .A1(opC13_out[17]), .A2(n3364), .Y(N1586) );
  AND2X1_RVT U1614 ( .A1(opC13_out[16]), .A2(n3364), .Y(N1585) );
  AND2X1_RVT U1615 ( .A1(opC13_out[15]), .A2(n3364), .Y(N1584) );
  AND2X1_RVT U1616 ( .A1(opC13_out[14]), .A2(n3364), .Y(N1583) );
  AND2X1_RVT U1617 ( .A1(opC13_out[13]), .A2(n3364), .Y(N1582) );
  AND2X1_RVT U1618 ( .A1(opC13_out[12]), .A2(n3364), .Y(N1581) );
  AND2X1_RVT U1619 ( .A1(opC13_out[11]), .A2(n3364), .Y(N1580) );
  AND2X1_RVT U1620 ( .A1(opC13_out[10]), .A2(n3364), .Y(N1579) );
  AND2X1_RVT U1621 ( .A1(opC13_out[9]), .A2(n3365), .Y(N1578) );
  AND2X1_RVT U1622 ( .A1(opC13_out[8]), .A2(n3365), .Y(N1577) );
  AND2X1_RVT U1623 ( .A1(opC13_out[7]), .A2(n3365), .Y(N1576) );
  AND2X1_RVT U1624 ( .A1(opC13_out[6]), .A2(n3365), .Y(N1575) );
  AND2X1_RVT U1625 ( .A1(opC13_out[5]), .A2(n3365), .Y(N1574) );
  AND2X1_RVT U1626 ( .A1(opC13_out[4]), .A2(n3365), .Y(N1573) );
  AND2X1_RVT U1627 ( .A1(opC13_out[3]), .A2(n3365), .Y(N1572) );
  AND2X1_RVT U1628 ( .A1(opC13_out[2]), .A2(n3365), .Y(N1571) );
  AND2X1_RVT U1629 ( .A1(opC13_out[1]), .A2(n3365), .Y(N1570) );
  AND2X1_RVT U1630 ( .A1(opC13_out[0]), .A2(n3365), .Y(N1569) );
  AND2X1_RVT U1631 ( .A1(opC30_out[31]), .A2(n3365), .Y(N1504) );
  AND2X1_RVT U1632 ( .A1(opC30_out[30]), .A2(n3365), .Y(N1503) );
  AND2X1_RVT U1633 ( .A1(opC30_out[29]), .A2(n3366), .Y(N1502) );
  AND2X1_RVT U1634 ( .A1(opC30_out[28]), .A2(n3366), .Y(N1501) );
  AND2X1_RVT U1635 ( .A1(opC30_out[27]), .A2(n3366), .Y(N1500) );
  AND2X1_RVT U1636 ( .A1(opC30_out[26]), .A2(n3366), .Y(N1499) );
  AND2X1_RVT U1637 ( .A1(opC30_out[25]), .A2(n3366), .Y(N1498) );
  AND2X1_RVT U1638 ( .A1(opC30_out[24]), .A2(n3366), .Y(N1497) );
  AND2X1_RVT U1639 ( .A1(opC30_out[23]), .A2(n3366), .Y(N1496) );
  AND2X1_RVT U1640 ( .A1(opC30_out[22]), .A2(n3366), .Y(N1495) );
  AND2X1_RVT U1641 ( .A1(opC30_out[21]), .A2(n3366), .Y(N1494) );
  AND2X1_RVT U1642 ( .A1(opC30_out[20]), .A2(n3366), .Y(N1493) );
  AND2X1_RVT U1643 ( .A1(opC30_out[19]), .A2(n3366), .Y(N1492) );
  AND2X1_RVT U1644 ( .A1(opC30_out[18]), .A2(n3366), .Y(N1491) );
  AND2X1_RVT U1645 ( .A1(opC30_out[17]), .A2(n3446), .Y(N1490) );
  AND2X1_RVT U1646 ( .A1(opC30_out[16]), .A2(n3447), .Y(N1489) );
  AND2X1_RVT U1647 ( .A1(opC30_out[15]), .A2(n3451), .Y(N1488) );
  AND2X1_RVT U1648 ( .A1(opC30_out[14]), .A2(n3452), .Y(N1487) );
  AND2X1_RVT U1649 ( .A1(opC30_out[13]), .A2(n3460), .Y(N1486) );
  AND2X1_RVT U1650 ( .A1(opC30_out[12]), .A2(n3448), .Y(N1485) );
  AND2X1_RVT U1651 ( .A1(opC30_out[11]), .A2(n3450), .Y(N1484) );
  AND2X1_RVT U1652 ( .A1(opC30_out[10]), .A2(n3449), .Y(N1483) );
  AND2X1_RVT U1653 ( .A1(opC30_out[9]), .A2(n3474), .Y(N1482) );
  AND2X1_RVT U1654 ( .A1(opC30_out[8]), .A2(n3453), .Y(N1481) );
  AND2X1_RVT U1655 ( .A1(opC30_out[7]), .A2(n3454), .Y(N1480) );
  AND2X1_RVT U1656 ( .A1(opC30_out[6]), .A2(n3466), .Y(N1479) );
  AND2X1_RVT U1657 ( .A1(opC30_out[5]), .A2(n3456), .Y(N1478) );
  AND2X1_RVT U1658 ( .A1(opC30_out[4]), .A2(n3458), .Y(N1477) );
  AND2X1_RVT U1659 ( .A1(opC30_out[3]), .A2(n3459), .Y(N1476) );
  AND2X1_RVT U1660 ( .A1(opC30_out[2]), .A2(n3460), .Y(N1475) );
  AND2X1_RVT U1661 ( .A1(opC30_out[1]), .A2(n3462), .Y(N1474) );
  AND2X1_RVT U1662 ( .A1(opC30_out[0]), .A2(n3474), .Y(N1473) );
  AND2X1_RVT U1663 ( .A1(opC21_out[31]), .A2(n3461), .Y(N1408) );
  AND2X1_RVT U1664 ( .A1(opC21_out[30]), .A2(n3463), .Y(N1407) );
  AND2X1_RVT U1665 ( .A1(opC21_out[29]), .A2(n3472), .Y(N1406) );
  AND2X1_RVT U1666 ( .A1(opC21_out[28]), .A2(n3442), .Y(N1405) );
  AND2X1_RVT U1667 ( .A1(opC21_out[27]), .A2(n3445), .Y(N1404) );
  AND2X1_RVT U1668 ( .A1(opC21_out[26]), .A2(n3466), .Y(N1403) );
  AND2X1_RVT U1669 ( .A1(opC21_out[25]), .A2(n3359), .Y(N1402) );
  AND2X1_RVT U1670 ( .A1(opC21_out[24]), .A2(n3364), .Y(N1401) );
  AND2X1_RVT U1671 ( .A1(opC21_out[23]), .A2(n3349), .Y(N1400) );
  AND2X1_RVT U1672 ( .A1(opC21_out[22]), .A2(n3349), .Y(N1399) );
  AND2X1_RVT U1673 ( .A1(opC21_out[21]), .A2(n3349), .Y(N1398) );
  AND2X1_RVT U1674 ( .A1(opC21_out[20]), .A2(n3349), .Y(N1397) );
  AND2X1_RVT U1675 ( .A1(opC21_out[19]), .A2(n3349), .Y(N1396) );
  AND2X1_RVT U1676 ( .A1(opC21_out[18]), .A2(n3349), .Y(N1395) );
  AND2X1_RVT U1677 ( .A1(opC21_out[17]), .A2(n3349), .Y(N1394) );
  AND2X1_RVT U1678 ( .A1(opC21_out[16]), .A2(n3349), .Y(N1393) );
  AND2X1_RVT U1679 ( .A1(opC21_out[15]), .A2(n3349), .Y(N1392) );
  AND2X1_RVT U1680 ( .A1(opC21_out[14]), .A2(n3349), .Y(N1391) );
  AND2X1_RVT U1681 ( .A1(opC21_out[13]), .A2(n3350), .Y(N1390) );
  AND2X1_RVT U1682 ( .A1(opC21_out[12]), .A2(n3350), .Y(N1389) );
  AND2X1_RVT U1683 ( .A1(opC21_out[11]), .A2(n3350), .Y(N1388) );
  AND2X1_RVT U1684 ( .A1(opC21_out[10]), .A2(n3350), .Y(N1387) );
  AND2X1_RVT U1685 ( .A1(opC21_out[9]), .A2(n3350), .Y(N1386) );
  AND2X1_RVT U1686 ( .A1(opC21_out[8]), .A2(n3466), .Y(N1385) );
  AND2X1_RVT U1687 ( .A1(opC21_out[7]), .A2(n3466), .Y(N1384) );
  AND2X1_RVT U1688 ( .A1(opC21_out[6]), .A2(n3466), .Y(N1383) );
  AND2X1_RVT U1689 ( .A1(opC21_out[5]), .A2(n3466), .Y(N1382) );
  AND2X1_RVT U1690 ( .A1(opC21_out[4]), .A2(n3466), .Y(N1381) );
  AND2X1_RVT U1691 ( .A1(opC21_out[3]), .A2(n3466), .Y(N1380) );
  AND2X1_RVT U1692 ( .A1(opC21_out[2]), .A2(n3466), .Y(N1379) );
  AND2X1_RVT U1693 ( .A1(opC21_out[1]), .A2(n3466), .Y(N1378) );
  AND2X1_RVT U1694 ( .A1(opC21_out[0]), .A2(n3466), .Y(N1377) );
  AND2X1_RVT U1695 ( .A1(opC12_out[31]), .A2(n3466), .Y(N1312) );
  AND2X1_RVT U1696 ( .A1(opC12_out[30]), .A2(n3466), .Y(N1311) );
  AND2X1_RVT U1697 ( .A1(opC12_out[29]), .A2(n3367), .Y(N1310) );
  AND2X1_RVT U1698 ( .A1(opC12_out[28]), .A2(n3367), .Y(N1309) );
  AND2X1_RVT U1699 ( .A1(opC12_out[27]), .A2(n3367), .Y(N1308) );
  AND2X1_RVT U1700 ( .A1(opC12_out[26]), .A2(n3367), .Y(N1307) );
  AND2X1_RVT U1701 ( .A1(opC12_out[25]), .A2(n3367), .Y(N1306) );
  AND2X1_RVT U1702 ( .A1(opC12_out[24]), .A2(n3369), .Y(N1305) );
  AND2X1_RVT U1703 ( .A1(opC12_out[23]), .A2(n3367), .Y(N1304) );
  AND2X1_RVT U1704 ( .A1(opC12_out[22]), .A2(n3367), .Y(N1303) );
  AND2X1_RVT U1705 ( .A1(opC12_out[21]), .A2(n3367), .Y(N1302) );
  AND2X1_RVT U1706 ( .A1(opC12_out[20]), .A2(n3367), .Y(N1301) );
  AND2X1_RVT U1707 ( .A1(opC12_out[19]), .A2(n3367), .Y(N1300) );
  AND2X1_RVT U1708 ( .A1(opC12_out[18]), .A2(n3367), .Y(N1299) );
  AND2X1_RVT U1709 ( .A1(opC12_out[17]), .A2(n3367), .Y(N1298) );
  AND2X1_RVT U1710 ( .A1(opC12_out[16]), .A2(n3347), .Y(N1297) );
  AND2X1_RVT U1711 ( .A1(opC12_out[15]), .A2(n3468), .Y(N1296) );
  AND2X1_RVT U1712 ( .A1(opC12_out[14]), .A2(n3368), .Y(N1295) );
  AND2X1_RVT U1713 ( .A1(opC12_out[13]), .A2(n3481), .Y(N1294) );
  AND2X1_RVT U1714 ( .A1(opC12_out[12]), .A2(n3442), .Y(N1293) );
  AND2X1_RVT U1715 ( .A1(opC12_out[11]), .A2(n3464), .Y(N1292) );
  AND2X1_RVT U1716 ( .A1(opC12_out[10]), .A2(n3480), .Y(N1291) );
  AND2X1_RVT U1717 ( .A1(opC12_out[9]), .A2(n3479), .Y(N1290) );
  AND2X1_RVT U1718 ( .A1(opC12_out[8]), .A2(n3477), .Y(N1289) );
  AND2X1_RVT U1719 ( .A1(opC12_out[7]), .A2(n3445), .Y(N1288) );
  AND2X1_RVT U1720 ( .A1(opC12_out[6]), .A2(n3443), .Y(N1287) );
  AND2X1_RVT U1721 ( .A1(opC12_out[5]), .A2(n3444), .Y(N1286) );
  AND2X1_RVT U1722 ( .A1(opC12_out[4]), .A2(n3368), .Y(N1285) );
  AND2X1_RVT U1723 ( .A1(opC12_out[3]), .A2(n3368), .Y(N1284) );
  AND2X1_RVT U1724 ( .A1(opC12_out[2]), .A2(n3368), .Y(N1283) );
  AND2X1_RVT U1725 ( .A1(opC12_out[1]), .A2(n3368), .Y(N1282) );
  AND2X1_RVT U1726 ( .A1(opC12_out[0]), .A2(n3368), .Y(N1281) );
  AND2X1_RVT U1727 ( .A1(opC03_out[31]), .A2(n3368), .Y(N1216) );
  AND2X1_RVT U1728 ( .A1(opC03_out[30]), .A2(n3368), .Y(N1215) );
  AND2X1_RVT U1729 ( .A1(opC03_out[29]), .A2(n3368), .Y(N1214) );
  AND2X1_RVT U1730 ( .A1(opC03_out[28]), .A2(n3368), .Y(N1213) );
  AND2X1_RVT U1731 ( .A1(opC03_out[27]), .A2(n3368), .Y(N1212) );
  AND2X1_RVT U1732 ( .A1(opC03_out[26]), .A2(n3368), .Y(N1211) );
  AND2X1_RVT U1733 ( .A1(opC03_out[25]), .A2(n3369), .Y(N1210) );
  AND2X1_RVT U1734 ( .A1(opC03_out[24]), .A2(n3369), .Y(N1209) );
  AND2X1_RVT U1735 ( .A1(opC03_out[23]), .A2(n3369), .Y(N1208) );
  AND2X1_RVT U1736 ( .A1(opC03_out[22]), .A2(n3369), .Y(N1207) );
  AND2X1_RVT U1737 ( .A1(opC03_out[21]), .A2(n3369), .Y(N1206) );
  AND2X1_RVT U1738 ( .A1(opC03_out[20]), .A2(n3369), .Y(N1205) );
  AND2X1_RVT U1739 ( .A1(opC03_out[19]), .A2(n3369), .Y(N1204) );
  AND2X1_RVT U1740 ( .A1(opC03_out[18]), .A2(n3369), .Y(N1203) );
  AND2X1_RVT U1741 ( .A1(opC03_out[17]), .A2(n3369), .Y(N1202) );
  AND2X1_RVT U1742 ( .A1(opC03_out[16]), .A2(n3369), .Y(N1201) );
  AND2X1_RVT U1743 ( .A1(opC03_out[15]), .A2(n3369), .Y(N1200) );
  AND2X1_RVT U1744 ( .A1(opC03_out[14]), .A2(n3370), .Y(N1199) );
  AND2X1_RVT U1745 ( .A1(opC03_out[13]), .A2(n3370), .Y(N1198) );
  AND2X1_RVT U1746 ( .A1(opC03_out[12]), .A2(n3370), .Y(N1197) );
  AND2X1_RVT U1747 ( .A1(opC03_out[11]), .A2(n3370), .Y(N1196) );
  AND2X1_RVT U1748 ( .A1(opC03_out[10]), .A2(n3370), .Y(N1195) );
  AND2X1_RVT U1749 ( .A1(opC03_out[9]), .A2(n3370), .Y(N1194) );
  AND2X1_RVT U1750 ( .A1(opC03_out[8]), .A2(n3370), .Y(N1193) );
  AND2X1_RVT U1751 ( .A1(opC03_out[7]), .A2(n3370), .Y(N1192) );
  AND2X1_RVT U1752 ( .A1(opC03_out[6]), .A2(n3370), .Y(N1191) );
  AND2X1_RVT U1753 ( .A1(opC03_out[5]), .A2(n3370), .Y(N1190) );
  AND2X1_RVT U1754 ( .A1(opC03_out[4]), .A2(n3370), .Y(N1189) );
  AND2X1_RVT U1755 ( .A1(opC03_out[3]), .A2(n3370), .Y(N1188) );
  AND2X1_RVT U1756 ( .A1(opC03_out[2]), .A2(n3371), .Y(N1187) );
  AND2X1_RVT U1757 ( .A1(opC03_out[1]), .A2(n3371), .Y(N1186) );
  AND2X1_RVT U1758 ( .A1(opC03_out[0]), .A2(n3371), .Y(N1185) );
  AND2X1_RVT U1759 ( .A1(opC20_out[31]), .A2(n3371), .Y(N1088) );
  AND2X1_RVT U1760 ( .A1(opC20_out[30]), .A2(n3371), .Y(N1087) );
  AND2X1_RVT U1761 ( .A1(opC20_out[29]), .A2(n3371), .Y(N1086) );
  AND2X1_RVT U1762 ( .A1(opC20_out[28]), .A2(n3371), .Y(N1085) );
  AND2X1_RVT U1763 ( .A1(opC20_out[27]), .A2(n3371), .Y(N1084) );
  AND2X1_RVT U1764 ( .A1(opC20_out[26]), .A2(n3371), .Y(N1083) );
  AND2X1_RVT U1765 ( .A1(opC20_out[25]), .A2(n3371), .Y(N1082) );
  AND2X1_RVT U1766 ( .A1(opC20_out[24]), .A2(n3371), .Y(N1081) );
  AND2X1_RVT U1767 ( .A1(opC20_out[23]), .A2(n3371), .Y(N1080) );
  AND2X1_RVT U1768 ( .A1(opC20_out[22]), .A2(n3464), .Y(N1079) );
  AND2X1_RVT U1769 ( .A1(opC20_out[21]), .A2(n3476), .Y(N1078) );
  AND2X1_RVT U1770 ( .A1(opC20_out[20]), .A2(n3457), .Y(N1077) );
  AND2X1_RVT U1771 ( .A1(opC20_out[19]), .A2(n3455), .Y(N1076) );
  AND2X1_RVT U1772 ( .A1(opC20_out[18]), .A2(n3481), .Y(N1075) );
  AND2X1_RVT U1773 ( .A1(opC20_out[17]), .A2(n3443), .Y(N1074) );
  AND2X1_RVT U1774 ( .A1(opC20_out[16]), .A2(n3444), .Y(N1073) );
  AND2X1_RVT U1775 ( .A1(opC20_out[15]), .A2(n3480), .Y(N1072) );
  AND2X1_RVT U1776 ( .A1(opC20_out[14]), .A2(n3478), .Y(N1071) );
  AND2X1_RVT U1777 ( .A1(opC20_out[13]), .A2(n3479), .Y(N1070) );
  AND2X1_RVT U1778 ( .A1(opC20_out[12]), .A2(n3477), .Y(N1069) );
  AND2X1_RVT U1779 ( .A1(opC20_out[11]), .A2(n3464), .Y(N1068) );
  AND2X1_RVT U1780 ( .A1(opC20_out[10]), .A2(n3474), .Y(N1067) );
  AND2X1_RVT U1781 ( .A1(opC20_out[9]), .A2(n3456), .Y(N1066) );
  AND2X1_RVT U1782 ( .A1(opC20_out[8]), .A2(n3458), .Y(N1065) );
  AND2X1_RVT U1783 ( .A1(opC20_out[7]), .A2(n3459), .Y(N1064) );
  AND2X1_RVT U1784 ( .A1(opC20_out[6]), .A2(n3460), .Y(N1063) );
  AND2X1_RVT U1785 ( .A1(opC20_out[5]), .A2(n3462), .Y(N1062) );
  AND2X1_RVT U1786 ( .A1(opC20_out[4]), .A2(n3461), .Y(N1061) );
  AND2X1_RVT U1787 ( .A1(opC20_out[3]), .A2(n3463), .Y(N1060) );
  AND2X1_RVT U1788 ( .A1(opC20_out[2]), .A2(n3441), .Y(N1059) );
  AND2X1_RVT U1789 ( .A1(opC20_out[1]), .A2(n3368), .Y(N1058) );
  AND2X1_RVT U1790 ( .A1(opC20_out[0]), .A2(n3466), .Y(N1057) );
  OSPEArray ospe_array ( .clk(clk), .rstnPipe(rstnPipe), .rstnPsum(rstnPsum), 
        .ipA0(ipA0), .ipA1(ipA1), .ipA2(ipA2), .ipA3(ipA3), .ipB0(ipB0), 
        .ipB1(ipB1), .ipB2(ipB2), .ipB3(ipB3), .opC00(opC00_out), .opC01(
        opC01_out), .opC02(opC02_out), .opC03(opC03_out), .opC10(opC10_out), 
        .opC11(opC11_out), .opC12(opC12_out), .opC13(opC13_out), .opC20(
        opC20_out), .opC21(opC21_out), .opC22(opC22_out), .opC23(opC23_out), 
        .opC30(opC30_out), .opC31(opC31_out), .opC32(opC32_out), .opC33(OpC33)
         );
  DATA_DW01_inc_0 add_46_S2 ( .A(BankAddr), .SUM({N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16}) );
  DFFX1_RVT opC00_d6_reg_31_ ( .D(n3215), .CLK(clk), .Q(n1073), .QN(n1074) );
  DFFX1_RVT opC00_d6_reg_30_ ( .D(n3214), .CLK(clk), .Q(n1072), .QN(n1075) );
  DFFX1_RVT opC00_d6_reg_29_ ( .D(n3213), .CLK(clk), .Q(n1071), .QN(n1076) );
  DFFX1_RVT opC00_d6_reg_28_ ( .D(n3212), .CLK(clk), .Q(n1070), .QN(n1077) );
  DFFX1_RVT opC00_d6_reg_27_ ( .D(n3211), .CLK(clk), .Q(n1069), .QN(n1078) );
  DFFX1_RVT opC00_d6_reg_26_ ( .D(n3210), .CLK(clk), .Q(n1068), .QN(n1079) );
  DFFX1_RVT opC00_d6_reg_25_ ( .D(n3209), .CLK(clk), .Q(n1067), .QN(n1080) );
  DFFX1_RVT opC00_d6_reg_24_ ( .D(n3208), .CLK(clk), .Q(n1066), .QN(n1081) );
  DFFX1_RVT opC00_d6_reg_23_ ( .D(n3207), .CLK(clk), .Q(n1065), .QN(n1082) );
  DFFX1_RVT opC00_d6_reg_22_ ( .D(n3206), .CLK(clk), .Q(n1064), .QN(n1083) );
  DFFX1_RVT opC00_d6_reg_21_ ( .D(n3205), .CLK(clk), .Q(n1063), .QN(n1084) );
  DFFX1_RVT opC00_d6_reg_20_ ( .D(n3204), .CLK(clk), .Q(n1062), .QN(n1085) );
  DFFX1_RVT opC00_d6_reg_19_ ( .D(n3203), .CLK(clk), .Q(n1061), .QN(n1086) );
  DFFX1_RVT opC00_d6_reg_18_ ( .D(n3202), .CLK(clk), .Q(n1060), .QN(n1087) );
  DFFX1_RVT opC00_d6_reg_17_ ( .D(n3201), .CLK(clk), .Q(n1059), .QN(n1088) );
  DFFX1_RVT opC00_d6_reg_16_ ( .D(n3200), .CLK(clk), .Q(n1058), .QN(n1089) );
  DFFX1_RVT opC00_d6_reg_15_ ( .D(n3199), .CLK(clk), .Q(n1057), .QN(n1090) );
  DFFX1_RVT opC00_d6_reg_14_ ( .D(n3198), .CLK(clk), .Q(n1056), .QN(n1091) );
  DFFX1_RVT opC00_d6_reg_13_ ( .D(n3197), .CLK(clk), .Q(n1055), .QN(n1092) );
  DFFX1_RVT opC00_d6_reg_12_ ( .D(n3196), .CLK(clk), .Q(n1054), .QN(n1093) );
  DFFX1_RVT opC00_d6_reg_11_ ( .D(n3195), .CLK(clk), .Q(n1053), .QN(n1094) );
  DFFX1_RVT opC00_d6_reg_10_ ( .D(n3194), .CLK(clk), .Q(n1052), .QN(n1095) );
  DFFX1_RVT opC00_d6_reg_9_ ( .D(n3193), .CLK(clk), .Q(n1051), .QN(n1096) );
  DFFX1_RVT opC00_d6_reg_8_ ( .D(n3192), .CLK(clk), .Q(n1050), .QN(n1097) );
  DFFX1_RVT opC00_d6_reg_7_ ( .D(n3191), .CLK(clk), .Q(n1049), .QN(n1098) );
  DFFX1_RVT opC00_d6_reg_6_ ( .D(n3190), .CLK(clk), .Q(n1048), .QN(n1099) );
  DFFX1_RVT opC00_d6_reg_5_ ( .D(n3189), .CLK(clk), .Q(n1047), .QN(n1100) );
  DFFX1_RVT opC00_d6_reg_4_ ( .D(n3188), .CLK(clk), .Q(n1046), .QN(n1101) );
  DFFX1_RVT opC00_d6_reg_3_ ( .D(n3187), .CLK(clk), .Q(n1045), .QN(n1102) );
  DFFX1_RVT opC00_d6_reg_2_ ( .D(n3186), .CLK(clk), .Q(n1044), .QN(n1103) );
  DFFX1_RVT opC00_d6_reg_1_ ( .D(n3185), .CLK(clk), .Q(n1043), .QN(n1104) );
  DFFX1_RVT opC00_d6_reg_0_ ( .D(n3184), .CLK(clk), .Q(n1042), .QN(n1105) );
  DFFX1_RVT BankAddr_reg_1_ ( .D(n3224), .CLK(clk), .Q(BankAddr[1]) );
  DFFX1_RVT BankAddr_reg_2_ ( .D(n3223), .CLK(clk), .Q(BankAddr[2]) );
  DFFX1_RVT BankAddr_reg_3_ ( .D(n3222), .CLK(clk), .Q(BankAddr[3]) );
  DFFX1_RVT BankAddr_reg_4_ ( .D(n3221), .CLK(clk), .Q(BankAddr[4]) );
  DFFX1_RVT BankAddr_reg_5_ ( .D(n3220), .CLK(clk), .Q(BankAddr[5]) );
  DFFX1_RVT BankAddr_reg_6_ ( .D(n3219), .CLK(clk), .Q(BankAddr[6]) );
  DFFX1_RVT BankAddr_reg_7_ ( .D(n3218), .CLK(clk), .Q(BankAddr[7]) );
  DFFX1_RVT BankAddr_reg_8_ ( .D(n3217), .CLK(clk), .Q(BankAddr[8]) );
  DFFX1_RVT BankAddr_reg_9_ ( .D(n3216), .CLK(clk), .Q(BankAddr[9]) );
  DFFX1_RVT BankAddr_reg_0_ ( .D(n3225), .CLK(clk), .Q(BankAddr[0]) );
  DFFX1_RVT opC01_d5_reg_31_ ( .D(N512), .CLK(clk), .QN(n2895) );
  DFFX1_RVT opC01_d5_reg_30_ ( .D(N511), .CLK(clk), .QN(n2894) );
  DFFX1_RVT opC01_d5_reg_29_ ( .D(N510), .CLK(clk), .QN(n2893) );
  DFFX1_RVT opC01_d5_reg_28_ ( .D(N509), .CLK(clk), .QN(n2892) );
  DFFX1_RVT opC01_d5_reg_27_ ( .D(N508), .CLK(clk), .QN(n2891) );
  DFFX1_RVT opC01_d5_reg_26_ ( .D(N507), .CLK(clk), .QN(n2890) );
  DFFX1_RVT opC01_d5_reg_25_ ( .D(N506), .CLK(clk), .QN(n2889) );
  DFFX1_RVT opC01_d5_reg_24_ ( .D(N505), .CLK(clk), .QN(n2888) );
  DFFX1_RVT opC01_d5_reg_23_ ( .D(N504), .CLK(clk), .QN(n2887) );
  DFFX1_RVT opC01_d5_reg_22_ ( .D(N503), .CLK(clk), .QN(n2886) );
  DFFX1_RVT opC01_d5_reg_21_ ( .D(N502), .CLK(clk), .QN(n2885) );
  DFFX1_RVT opC01_d5_reg_20_ ( .D(N501), .CLK(clk), .QN(n2884) );
  DFFX1_RVT opC01_d5_reg_19_ ( .D(N500), .CLK(clk), .QN(n2883) );
  DFFX1_RVT opC01_d5_reg_18_ ( .D(N499), .CLK(clk), .QN(n2882) );
  DFFX1_RVT opC01_d5_reg_17_ ( .D(N498), .CLK(clk), .QN(n2881) );
  DFFX1_RVT opC01_d5_reg_16_ ( .D(N497), .CLK(clk), .QN(n2880) );
  DFFX1_RVT opC01_d5_reg_15_ ( .D(N496), .CLK(clk), .QN(n2879) );
  DFFX1_RVT opC01_d5_reg_14_ ( .D(N495), .CLK(clk), .QN(n2878) );
  DFFX1_RVT opC01_d5_reg_13_ ( .D(N494), .CLK(clk), .QN(n2877) );
  DFFX1_RVT opC01_d5_reg_12_ ( .D(N493), .CLK(clk), .QN(n2876) );
  DFFX1_RVT opC01_d5_reg_11_ ( .D(N492), .CLK(clk), .QN(n2875) );
  DFFX1_RVT opC01_d5_reg_10_ ( .D(N491), .CLK(clk), .QN(n2874) );
  DFFX1_RVT opC01_d5_reg_9_ ( .D(N490), .CLK(clk), .QN(n2873) );
  DFFX1_RVT opC01_d5_reg_8_ ( .D(N489), .CLK(clk), .QN(n2872) );
  DFFX1_RVT opC01_d5_reg_7_ ( .D(N488), .CLK(clk), .QN(n2871) );
  DFFX1_RVT opC01_d5_reg_6_ ( .D(N487), .CLK(clk), .QN(n2870) );
  DFFX1_RVT opC01_d5_reg_5_ ( .D(N486), .CLK(clk), .QN(n2869) );
  DFFX1_RVT opC01_d5_reg_4_ ( .D(N485), .CLK(clk), .QN(n2868) );
  DFFX1_RVT opC01_d5_reg_3_ ( .D(N484), .CLK(clk), .QN(n2867) );
  DFFX1_RVT opC01_d5_reg_2_ ( .D(N483), .CLK(clk), .QN(n2866) );
  DFFX1_RVT opC01_d5_reg_1_ ( .D(N482), .CLK(clk), .QN(n2865) );
  DFFX1_RVT opC01_d5_reg_0_ ( .D(N481), .CLK(clk), .QN(n2864) );
  DFFX1_RVT opC10_d5_reg_31_ ( .D(N672), .CLK(clk), .QN(n2639) );
  DFFX1_RVT opC10_d5_reg_30_ ( .D(N671), .CLK(clk), .QN(n2638) );
  DFFX1_RVT opC10_d5_reg_29_ ( .D(N670), .CLK(clk), .QN(n2637) );
  DFFX1_RVT opC10_d5_reg_28_ ( .D(N669), .CLK(clk), .QN(n2636) );
  DFFX1_RVT opC10_d5_reg_27_ ( .D(N668), .CLK(clk), .QN(n2635) );
  DFFX1_RVT opC10_d5_reg_26_ ( .D(N667), .CLK(clk), .QN(n2634) );
  DFFX1_RVT opC10_d5_reg_25_ ( .D(N666), .CLK(clk), .QN(n2633) );
  DFFX1_RVT opC10_d5_reg_24_ ( .D(N665), .CLK(clk), .QN(n2632) );
  DFFX1_RVT opC10_d5_reg_23_ ( .D(N664), .CLK(clk), .QN(n2631) );
  DFFX1_RVT opC10_d5_reg_22_ ( .D(N663), .CLK(clk), .QN(n2630) );
  DFFX1_RVT opC10_d5_reg_21_ ( .D(N662), .CLK(clk), .QN(n2629) );
  DFFX1_RVT opC10_d5_reg_20_ ( .D(N661), .CLK(clk), .QN(n2628) );
  DFFX1_RVT opC10_d5_reg_19_ ( .D(N660), .CLK(clk), .QN(n2627) );
  DFFX1_RVT opC10_d5_reg_18_ ( .D(N659), .CLK(clk), .QN(n2626) );
  DFFX1_RVT opC10_d5_reg_17_ ( .D(N658), .CLK(clk), .QN(n2625) );
  DFFX1_RVT opC10_d5_reg_16_ ( .D(N657), .CLK(clk), .QN(n2624) );
  DFFX1_RVT opC10_d5_reg_15_ ( .D(N656), .CLK(clk), .QN(n2623) );
  DFFX1_RVT opC10_d5_reg_14_ ( .D(N655), .CLK(clk), .QN(n2622) );
  DFFX1_RVT opC10_d5_reg_13_ ( .D(N654), .CLK(clk), .QN(n2621) );
  DFFX1_RVT opC10_d5_reg_12_ ( .D(N653), .CLK(clk), .QN(n2620) );
  DFFX1_RVT opC10_d5_reg_11_ ( .D(N652), .CLK(clk), .QN(n2619) );
  DFFX1_RVT opC10_d5_reg_10_ ( .D(N651), .CLK(clk), .QN(n2618) );
  DFFX1_RVT opC10_d5_reg_9_ ( .D(N650), .CLK(clk), .QN(n2617) );
  DFFX1_RVT opC10_d5_reg_8_ ( .D(N649), .CLK(clk), .QN(n2616) );
  DFFX1_RVT opC10_d5_reg_7_ ( .D(N648), .CLK(clk), .QN(n2615) );
  DFFX1_RVT opC10_d5_reg_6_ ( .D(N647), .CLK(clk), .QN(n2614) );
  DFFX1_RVT opC10_d5_reg_5_ ( .D(N646), .CLK(clk), .QN(n2613) );
  DFFX1_RVT opC10_d5_reg_4_ ( .D(N645), .CLK(clk), .QN(n2612) );
  DFFX1_RVT opC10_d5_reg_3_ ( .D(N644), .CLK(clk), .QN(n2611) );
  DFFX1_RVT opC10_d5_reg_2_ ( .D(N643), .CLK(clk), .QN(n2610) );
  DFFX1_RVT opC10_d5_reg_1_ ( .D(N642), .CLK(clk), .QN(n2609) );
  DFFX1_RVT opC10_d5_reg_0_ ( .D(N641), .CLK(clk), .QN(n2608) );
  DFFX1_RVT opC02_d4_reg_31_ ( .D(N832), .CLK(clk), .QN(n2383) );
  DFFX1_RVT opC02_d4_reg_30_ ( .D(N831), .CLK(clk), .QN(n2382) );
  DFFX1_RVT opC02_d4_reg_29_ ( .D(N830), .CLK(clk), .QN(n2381) );
  DFFX1_RVT opC02_d4_reg_28_ ( .D(N829), .CLK(clk), .QN(n2380) );
  DFFX1_RVT opC02_d4_reg_27_ ( .D(N828), .CLK(clk), .QN(n2379) );
  DFFX1_RVT opC02_d4_reg_26_ ( .D(N827), .CLK(clk), .QN(n2378) );
  DFFX1_RVT opC02_d4_reg_25_ ( .D(N826), .CLK(clk), .QN(n2377) );
  DFFX1_RVT opC02_d4_reg_24_ ( .D(N825), .CLK(clk), .QN(n2376) );
  DFFX1_RVT opC02_d4_reg_23_ ( .D(N824), .CLK(clk), .QN(n2375) );
  DFFX1_RVT opC02_d4_reg_22_ ( .D(N823), .CLK(clk), .QN(n2374) );
  DFFX1_RVT opC02_d4_reg_21_ ( .D(N822), .CLK(clk), .QN(n2373) );
  DFFX1_RVT opC02_d4_reg_20_ ( .D(N821), .CLK(clk), .QN(n2372) );
  DFFX1_RVT opC02_d4_reg_19_ ( .D(N820), .CLK(clk), .QN(n2371) );
  DFFX1_RVT opC02_d4_reg_18_ ( .D(N819), .CLK(clk), .QN(n2370) );
  DFFX1_RVT opC02_d4_reg_17_ ( .D(N818), .CLK(clk), .QN(n2369) );
  DFFX1_RVT opC02_d4_reg_16_ ( .D(N817), .CLK(clk), .QN(n2368) );
  DFFX1_RVT opC02_d4_reg_15_ ( .D(N816), .CLK(clk), .QN(n2367) );
  DFFX1_RVT opC02_d4_reg_14_ ( .D(N815), .CLK(clk), .QN(n2366) );
  DFFX1_RVT opC02_d4_reg_13_ ( .D(N814), .CLK(clk), .QN(n2365) );
  DFFX1_RVT opC02_d4_reg_12_ ( .D(N813), .CLK(clk), .QN(n2364) );
  DFFX1_RVT opC02_d4_reg_11_ ( .D(N812), .CLK(clk), .QN(n2363) );
  DFFX1_RVT opC02_d4_reg_10_ ( .D(N811), .CLK(clk), .QN(n2362) );
  DFFX1_RVT opC02_d4_reg_9_ ( .D(N810), .CLK(clk), .QN(n2361) );
  DFFX1_RVT opC02_d4_reg_8_ ( .D(N809), .CLK(clk), .QN(n2360) );
  DFFX1_RVT opC02_d4_reg_7_ ( .D(N808), .CLK(clk), .QN(n2359) );
  DFFX1_RVT opC02_d4_reg_6_ ( .D(N807), .CLK(clk), .QN(n2358) );
  DFFX1_RVT opC02_d4_reg_5_ ( .D(N806), .CLK(clk), .QN(n2357) );
  DFFX1_RVT opC02_d4_reg_4_ ( .D(N805), .CLK(clk), .QN(n2356) );
  DFFX1_RVT opC02_d4_reg_3_ ( .D(N804), .CLK(clk), .QN(n2355) );
  DFFX1_RVT opC02_d4_reg_2_ ( .D(N803), .CLK(clk), .QN(n2354) );
  DFFX1_RVT opC02_d4_reg_1_ ( .D(N802), .CLK(clk), .QN(n2353) );
  DFFX1_RVT opC02_d4_reg_0_ ( .D(N801), .CLK(clk), .QN(n2352) );
  DFFX1_RVT opC11_d4_reg_31_ ( .D(N960), .CLK(clk), .QN(n2191) );
  DFFX1_RVT opC11_d4_reg_30_ ( .D(N959), .CLK(clk), .QN(n2190) );
  DFFX1_RVT opC11_d4_reg_29_ ( .D(N958), .CLK(clk), .QN(n2189) );
  DFFX1_RVT opC11_d4_reg_28_ ( .D(N957), .CLK(clk), .QN(n2188) );
  DFFX1_RVT opC11_d4_reg_27_ ( .D(N956), .CLK(clk), .QN(n2187) );
  DFFX1_RVT opC11_d4_reg_26_ ( .D(N955), .CLK(clk), .QN(n2186) );
  DFFX1_RVT opC11_d4_reg_25_ ( .D(N954), .CLK(clk), .QN(n2185) );
  DFFX1_RVT opC11_d4_reg_24_ ( .D(N953), .CLK(clk), .QN(n2184) );
  DFFX1_RVT opC11_d4_reg_23_ ( .D(N952), .CLK(clk), .QN(n2183) );
  DFFX1_RVT opC11_d4_reg_22_ ( .D(N951), .CLK(clk), .QN(n2182) );
  DFFX1_RVT opC11_d4_reg_21_ ( .D(N950), .CLK(clk), .QN(n2181) );
  DFFX1_RVT opC11_d4_reg_20_ ( .D(N949), .CLK(clk), .QN(n2180) );
  DFFX1_RVT opC11_d4_reg_19_ ( .D(N948), .CLK(clk), .QN(n2179) );
  DFFX1_RVT opC11_d4_reg_18_ ( .D(N947), .CLK(clk), .QN(n2178) );
  DFFX1_RVT opC11_d4_reg_17_ ( .D(N946), .CLK(clk), .QN(n2177) );
  DFFX1_RVT opC11_d4_reg_16_ ( .D(N945), .CLK(clk), .QN(n2176) );
  DFFX1_RVT opC11_d4_reg_15_ ( .D(N944), .CLK(clk), .QN(n2175) );
  DFFX1_RVT opC11_d4_reg_14_ ( .D(N943), .CLK(clk), .QN(n2174) );
  DFFX1_RVT opC11_d4_reg_13_ ( .D(N942), .CLK(clk), .QN(n2173) );
  DFFX1_RVT opC11_d4_reg_12_ ( .D(N941), .CLK(clk), .QN(n2172) );
  DFFX1_RVT opC11_d4_reg_11_ ( .D(N940), .CLK(clk), .QN(n2171) );
  DFFX1_RVT opC11_d4_reg_10_ ( .D(N939), .CLK(clk), .QN(n2170) );
  DFFX1_RVT opC11_d4_reg_9_ ( .D(N938), .CLK(clk), .QN(n2169) );
  DFFX1_RVT opC11_d4_reg_8_ ( .D(N937), .CLK(clk), .QN(n2168) );
  DFFX1_RVT opC11_d4_reg_7_ ( .D(N936), .CLK(clk), .QN(n2167) );
  DFFX1_RVT opC11_d4_reg_6_ ( .D(N935), .CLK(clk), .QN(n2166) );
  DFFX1_RVT opC11_d4_reg_5_ ( .D(N934), .CLK(clk), .QN(n2165) );
  DFFX1_RVT opC11_d4_reg_4_ ( .D(N933), .CLK(clk), .QN(n2164) );
  DFFX1_RVT opC11_d4_reg_3_ ( .D(N932), .CLK(clk), .QN(n2163) );
  DFFX1_RVT opC11_d4_reg_2_ ( .D(N931), .CLK(clk), .QN(n2162) );
  DFFX1_RVT opC11_d4_reg_1_ ( .D(N930), .CLK(clk), .QN(n2161) );
  DFFX1_RVT opC11_d2_reg_6_ ( .D(N999), .CLK(clk), .QN(n2046) );
  DFFX1_RVT opC20_d4_reg_31_ ( .D(N1088), .CLK(clk), .QN(n2001) );
  DFFX1_RVT opC20_d4_reg_30_ ( .D(N1087), .CLK(clk), .QN(n2000) );
  DFFX1_RVT opC20_d4_reg_29_ ( .D(N1086), .CLK(clk), .QN(n1999) );
  DFFX1_RVT opC20_d4_reg_28_ ( .D(N1085), .CLK(clk), .QN(n1998) );
  DFFX1_RVT opC20_d4_reg_27_ ( .D(N1084), .CLK(clk), .QN(n1997) );
  DFFX1_RVT opC20_d4_reg_26_ ( .D(N1083), .CLK(clk), .QN(n1996) );
  DFFX1_RVT opC20_d4_reg_25_ ( .D(N1082), .CLK(clk), .QN(n1995) );
  DFFX1_RVT opC20_d4_reg_24_ ( .D(N1081), .CLK(clk), .QN(n1994) );
  DFFX1_RVT opC20_d4_reg_23_ ( .D(N1080), .CLK(clk), .QN(n1993) );
  DFFX1_RVT opC20_d4_reg_22_ ( .D(N1079), .CLK(clk), .QN(n1992) );
  DFFX1_RVT opC20_d4_reg_21_ ( .D(N1078), .CLK(clk), .QN(n1991) );
  DFFX1_RVT opC20_d4_reg_20_ ( .D(N1077), .CLK(clk), .QN(n1990) );
  DFFX1_RVT opC20_d4_reg_19_ ( .D(N1076), .CLK(clk), .QN(n1989) );
  DFFX1_RVT opC20_d4_reg_18_ ( .D(N1075), .CLK(clk), .QN(n1988) );
  DFFX1_RVT opC20_d4_reg_17_ ( .D(N1074), .CLK(clk), .QN(n1987) );
  DFFX1_RVT opC20_d4_reg_16_ ( .D(N1073), .CLK(clk), .QN(n1986) );
  DFFX1_RVT opC20_d4_reg_15_ ( .D(N1072), .CLK(clk), .QN(n1985) );
  DFFX1_RVT opC20_d4_reg_14_ ( .D(N1071), .CLK(clk), .QN(n1984) );
  DFFX1_RVT opC20_d4_reg_13_ ( .D(N1070), .CLK(clk), .QN(n1983) );
  DFFX1_RVT opC20_d4_reg_12_ ( .D(N1069), .CLK(clk), .QN(n1982) );
  DFFX1_RVT opC20_d4_reg_11_ ( .D(N1068), .CLK(clk), .QN(n1981) );
  DFFX1_RVT opC20_d4_reg_10_ ( .D(N1067), .CLK(clk), .QN(n1980) );
  DFFX1_RVT opC20_d4_reg_9_ ( .D(N1066), .CLK(clk), .QN(n1979) );
  DFFX1_RVT opC20_d4_reg_8_ ( .D(N1065), .CLK(clk), .QN(n1978) );
  DFFX1_RVT opC20_d4_reg_7_ ( .D(N1064), .CLK(clk), .QN(n1977) );
  DFFX1_RVT opC20_d4_reg_6_ ( .D(N1063), .CLK(clk), .QN(n1976) );
  DFFX1_RVT opC20_d4_reg_5_ ( .D(N1062), .CLK(clk), .QN(n1975) );
  DFFX1_RVT opC20_d4_reg_4_ ( .D(N1061), .CLK(clk), .QN(n1974) );
  DFFX1_RVT opC20_d4_reg_3_ ( .D(N1060), .CLK(clk), .QN(n1973) );
  DFFX1_RVT opC20_d4_reg_2_ ( .D(N1059), .CLK(clk), .QN(n1972) );
  DFFX1_RVT opC20_d4_reg_1_ ( .D(N1058), .CLK(clk), .QN(n1971) );
  DFFX1_RVT opC20_d4_reg_0_ ( .D(N1057), .CLK(clk), .QN(n1970) );
  DFFX1_RVT opC03_d3_reg_31_ ( .D(N1216), .CLK(clk), .QN(n1809) );
  DFFX1_RVT opC03_d3_reg_30_ ( .D(N1215), .CLK(clk), .QN(n1808) );
  DFFX1_RVT opC03_d3_reg_29_ ( .D(N1214), .CLK(clk), .QN(n1807) );
  DFFX1_RVT opC03_d3_reg_28_ ( .D(N1213), .CLK(clk), .QN(n1806) );
  DFFX1_RVT opC03_d3_reg_27_ ( .D(N1212), .CLK(clk), .QN(n1805) );
  DFFX1_RVT opC03_d3_reg_26_ ( .D(N1211), .CLK(clk), .QN(n1804) );
  DFFX1_RVT opC03_d3_reg_25_ ( .D(N1210), .CLK(clk), .QN(n1803) );
  DFFX1_RVT opC03_d3_reg_24_ ( .D(N1209), .CLK(clk), .QN(n1802) );
  DFFX1_RVT opC03_d3_reg_23_ ( .D(N1208), .CLK(clk), .QN(n1801) );
  DFFX1_RVT opC03_d3_reg_22_ ( .D(N1207), .CLK(clk), .QN(n1800) );
  DFFX1_RVT opC03_d3_reg_21_ ( .D(N1206), .CLK(clk), .QN(n1799) );
  DFFX1_RVT opC03_d3_reg_20_ ( .D(N1205), .CLK(clk), .QN(n1798) );
  DFFX1_RVT opC03_d3_reg_19_ ( .D(N1204), .CLK(clk), .QN(n1797) );
  DFFX1_RVT opC03_d3_reg_18_ ( .D(N1203), .CLK(clk), .QN(n1796) );
  DFFX1_RVT opC03_d3_reg_17_ ( .D(N1202), .CLK(clk), .QN(n1795) );
  DFFX1_RVT opC03_d3_reg_16_ ( .D(N1201), .CLK(clk), .QN(n1794) );
  DFFX1_RVT opC03_d3_reg_15_ ( .D(N1200), .CLK(clk), .QN(n1793) );
  DFFX1_RVT opC03_d3_reg_14_ ( .D(N1199), .CLK(clk), .QN(n1792) );
  DFFX1_RVT opC03_d3_reg_13_ ( .D(N1198), .CLK(clk), .QN(n1791) );
  DFFX1_RVT opC03_d3_reg_12_ ( .D(N1197), .CLK(clk), .QN(n1790) );
  DFFX1_RVT opC03_d3_reg_11_ ( .D(N1196), .CLK(clk), .QN(n1789) );
  DFFX1_RVT opC03_d3_reg_10_ ( .D(N1195), .CLK(clk), .QN(n1788) );
  DFFX1_RVT opC03_d3_reg_9_ ( .D(N1194), .CLK(clk), .QN(n1787) );
  DFFX1_RVT opC03_d3_reg_8_ ( .D(N1193), .CLK(clk), .QN(n1786) );
  DFFX1_RVT opC03_d3_reg_7_ ( .D(N1192), .CLK(clk), .QN(n1785) );
  DFFX1_RVT opC03_d3_reg_6_ ( .D(N1191), .CLK(clk), .QN(n1784) );
  DFFX1_RVT opC03_d3_reg_5_ ( .D(N1190), .CLK(clk), .QN(n1783) );
  DFFX1_RVT opC03_d3_reg_4_ ( .D(N1189), .CLK(clk), .QN(n1782) );
  DFFX1_RVT opC03_d3_reg_3_ ( .D(N1188), .CLK(clk), .QN(n1781) );
  DFFX1_RVT opC03_d3_reg_2_ ( .D(N1187), .CLK(clk), .QN(n1780) );
  DFFX1_RVT opC03_d3_reg_1_ ( .D(N1186), .CLK(clk), .QN(n1779) );
  DFFX1_RVT opC03_d3_reg_0_ ( .D(N1185), .CLK(clk), .QN(n1778) );
  DFFX1_RVT opC12_d3_reg_31_ ( .D(N1312), .CLK(clk), .QN(n1681) );
  DFFX1_RVT opC12_d3_reg_30_ ( .D(N1311), .CLK(clk), .QN(n1680) );
  DFFX1_RVT opC12_d3_reg_29_ ( .D(N1310), .CLK(clk), .QN(n1679) );
  DFFX1_RVT opC12_d3_reg_28_ ( .D(N1309), .CLK(clk), .QN(n1678) );
  DFFX1_RVT opC12_d3_reg_27_ ( .D(N1308), .CLK(clk), .QN(n1677) );
  DFFX1_RVT opC12_d3_reg_26_ ( .D(N1307), .CLK(clk), .QN(n1676) );
  DFFX1_RVT opC12_d3_reg_25_ ( .D(N1306), .CLK(clk), .QN(n1675) );
  DFFX1_RVT opC12_d3_reg_24_ ( .D(N1305), .CLK(clk), .QN(n1674) );
  DFFX1_RVT opC12_d3_reg_23_ ( .D(N1304), .CLK(clk), .QN(n1673) );
  DFFX1_RVT opC12_d3_reg_22_ ( .D(N1303), .CLK(clk), .QN(n1672) );
  DFFX1_RVT opC12_d3_reg_21_ ( .D(N1302), .CLK(clk), .QN(n1671) );
  DFFX1_RVT opC12_d3_reg_20_ ( .D(N1301), .CLK(clk), .QN(n1670) );
  DFFX1_RVT opC12_d3_reg_19_ ( .D(N1300), .CLK(clk), .QN(n1669) );
  DFFX1_RVT opC12_d3_reg_18_ ( .D(N1299), .CLK(clk), .QN(n1668) );
  DFFX1_RVT opC12_d3_reg_17_ ( .D(N1298), .CLK(clk), .QN(n1667) );
  DFFX1_RVT opC12_d3_reg_16_ ( .D(N1297), .CLK(clk), .QN(n1666) );
  DFFX1_RVT opC12_d3_reg_15_ ( .D(N1296), .CLK(clk), .QN(n1665) );
  DFFX1_RVT opC12_d3_reg_14_ ( .D(N1295), .CLK(clk), .QN(n1664) );
  DFFX1_RVT opC12_d3_reg_13_ ( .D(N1294), .CLK(clk), .QN(n1663) );
  DFFX1_RVT opC12_d3_reg_12_ ( .D(N1293), .CLK(clk), .QN(n1662) );
  DFFX1_RVT opC12_d3_reg_11_ ( .D(N1292), .CLK(clk), .QN(n1661) );
  DFFX1_RVT opC12_d3_reg_10_ ( .D(N1291), .CLK(clk), .QN(n1660) );
  DFFX1_RVT opC12_d3_reg_9_ ( .D(N1290), .CLK(clk), .QN(n1659) );
  DFFX1_RVT opC12_d3_reg_8_ ( .D(N1289), .CLK(clk), .QN(n1658) );
  DFFX1_RVT opC12_d3_reg_7_ ( .D(N1288), .CLK(clk), .QN(n1657) );
  DFFX1_RVT opC12_d3_reg_6_ ( .D(N1287), .CLK(clk), .QN(n1656) );
  DFFX1_RVT opC12_d3_reg_5_ ( .D(N1286), .CLK(clk), .QN(n1655) );
  DFFX1_RVT opC12_d3_reg_4_ ( .D(N1285), .CLK(clk), .QN(n1654) );
  DFFX1_RVT opC12_d3_reg_3_ ( .D(N1284), .CLK(clk), .QN(n1653) );
  DFFX1_RVT opC12_d3_reg_2_ ( .D(N1283), .CLK(clk), .QN(n1652) );
  DFFX1_RVT opC12_d3_reg_1_ ( .D(N1282), .CLK(clk), .QN(n1651) );
  DFFX1_RVT opC12_d3_reg_0_ ( .D(N1281), .CLK(clk), .QN(n1650) );
  DFFX1_RVT opC21_d3_reg_31_ ( .D(N1408), .CLK(clk), .QN(n1553) );
  DFFX1_RVT opC21_d3_reg_30_ ( .D(N1407), .CLK(clk), .QN(n1552) );
  DFFX1_RVT opC21_d3_reg_29_ ( .D(N1406), .CLK(clk), .QN(n1551) );
  DFFX1_RVT opC21_d3_reg_28_ ( .D(N1405), .CLK(clk), .QN(n1550) );
  DFFX1_RVT opC21_d3_reg_27_ ( .D(N1404), .CLK(clk), .QN(n1549) );
  DFFX1_RVT opC21_d3_reg_26_ ( .D(N1403), .CLK(clk), .QN(n1548) );
  DFFX1_RVT opC21_d3_reg_25_ ( .D(N1402), .CLK(clk), .QN(n1547) );
  DFFX1_RVT opC21_d3_reg_24_ ( .D(N1401), .CLK(clk), .QN(n1546) );
  DFFX1_RVT opC21_d3_reg_23_ ( .D(N1400), .CLK(clk), .QN(n1545) );
  DFFX1_RVT opC21_d3_reg_22_ ( .D(N1399), .CLK(clk), .QN(n1544) );
  DFFX1_RVT opC21_d3_reg_21_ ( .D(N1398), .CLK(clk), .QN(n1543) );
  DFFX1_RVT opC21_d3_reg_20_ ( .D(N1397), .CLK(clk), .QN(n1542) );
  DFFX1_RVT opC21_d3_reg_19_ ( .D(N1396), .CLK(clk), .QN(n1541) );
  DFFX1_RVT opC21_d3_reg_18_ ( .D(N1395), .CLK(clk), .QN(n1540) );
  DFFX1_RVT opC21_d3_reg_17_ ( .D(N1394), .CLK(clk), .QN(n1539) );
  DFFX1_RVT opC21_d3_reg_16_ ( .D(N1393), .CLK(clk), .QN(n1538) );
  DFFX1_RVT opC21_d3_reg_15_ ( .D(N1392), .CLK(clk), .QN(n1537) );
  DFFX1_RVT opC21_d3_reg_14_ ( .D(N1391), .CLK(clk), .QN(n1536) );
  DFFX1_RVT opC21_d3_reg_13_ ( .D(N1390), .CLK(clk), .QN(n1535) );
  DFFX1_RVT opC21_d3_reg_12_ ( .D(N1389), .CLK(clk), .QN(n1534) );
  DFFX1_RVT opC21_d3_reg_11_ ( .D(N1388), .CLK(clk), .QN(n1533) );
  DFFX1_RVT opC21_d3_reg_10_ ( .D(N1387), .CLK(clk), .QN(n1532) );
  DFFX1_RVT opC21_d3_reg_9_ ( .D(N1386), .CLK(clk), .QN(n1531) );
  DFFX1_RVT opC21_d3_reg_8_ ( .D(N1385), .CLK(clk), .QN(n1530) );
  DFFX1_RVT opC21_d3_reg_7_ ( .D(N1384), .CLK(clk), .QN(n1529) );
  DFFX1_RVT opC21_d3_reg_6_ ( .D(N1383), .CLK(clk), .QN(n1528) );
  DFFX1_RVT opC21_d3_reg_5_ ( .D(N1382), .CLK(clk), .QN(n1527) );
  DFFX1_RVT opC21_d3_reg_4_ ( .D(N1381), .CLK(clk), .QN(n1526) );
  DFFX1_RVT opC21_d3_reg_3_ ( .D(N1380), .CLK(clk), .QN(n1525) );
  DFFX1_RVT opC21_d3_reg_2_ ( .D(N1379), .CLK(clk), .QN(n1524) );
  DFFX1_RVT opC21_d3_reg_1_ ( .D(N1378), .CLK(clk), .QN(n1523) );
  DFFX1_RVT opC21_d3_reg_0_ ( .D(N1377), .CLK(clk), .QN(n1522) );
  DFFX1_RVT opC30_d3_reg_31_ ( .D(N1504), .CLK(clk), .QN(n1425) );
  DFFX1_RVT opC30_d3_reg_30_ ( .D(N1503), .CLK(clk), .QN(n1424) );
  DFFX1_RVT opC30_d3_reg_29_ ( .D(N1502), .CLK(clk), .QN(n1423) );
  DFFX1_RVT opC30_d3_reg_28_ ( .D(N1501), .CLK(clk), .QN(n1422) );
  DFFX1_RVT opC30_d3_reg_27_ ( .D(N1500), .CLK(clk), .QN(n1421) );
  DFFX1_RVT opC30_d3_reg_26_ ( .D(N1499), .CLK(clk), .QN(n1420) );
  DFFX1_RVT opC30_d3_reg_25_ ( .D(N1498), .CLK(clk), .QN(n1419) );
  DFFX1_RVT opC30_d3_reg_24_ ( .D(N1497), .CLK(clk), .QN(n1418) );
  DFFX1_RVT opC30_d3_reg_23_ ( .D(N1496), .CLK(clk), .QN(n1417) );
  DFFX1_RVT opC30_d3_reg_22_ ( .D(N1495), .CLK(clk), .QN(n1416) );
  DFFX1_RVT opC30_d3_reg_21_ ( .D(N1494), .CLK(clk), .QN(n1415) );
  DFFX1_RVT opC30_d3_reg_20_ ( .D(N1493), .CLK(clk), .QN(n1414) );
  DFFX1_RVT opC30_d3_reg_19_ ( .D(N1492), .CLK(clk), .QN(n1413) );
  DFFX1_RVT opC30_d3_reg_18_ ( .D(N1491), .CLK(clk), .QN(n1412) );
  DFFX1_RVT opC30_d3_reg_17_ ( .D(N1490), .CLK(clk), .QN(n1411) );
  DFFX1_RVT opC30_d3_reg_16_ ( .D(N1489), .CLK(clk), .QN(n1410) );
  DFFX1_RVT opC30_d3_reg_15_ ( .D(N1488), .CLK(clk), .QN(n1409) );
  DFFX1_RVT opC30_d3_reg_14_ ( .D(N1487), .CLK(clk), .QN(n1408) );
  DFFX1_RVT opC30_d3_reg_13_ ( .D(N1486), .CLK(clk), .QN(n1407) );
  DFFX1_RVT opC30_d3_reg_12_ ( .D(N1485), .CLK(clk), .QN(n1406) );
  DFFX1_RVT opC30_d3_reg_11_ ( .D(N1484), .CLK(clk), .QN(n1405) );
  DFFX1_RVT opC30_d3_reg_10_ ( .D(N1483), .CLK(clk), .QN(n1404) );
  DFFX1_RVT opC30_d3_reg_9_ ( .D(N1482), .CLK(clk), .QN(n1403) );
  DFFX1_RVT opC30_d3_reg_8_ ( .D(N1481), .CLK(clk), .QN(n1402) );
  DFFX1_RVT opC30_d3_reg_7_ ( .D(N1480), .CLK(clk), .QN(n1401) );
  DFFX1_RVT opC30_d3_reg_6_ ( .D(N1479), .CLK(clk), .QN(n1400) );
  DFFX1_RVT opC30_d3_reg_5_ ( .D(N1478), .CLK(clk), .QN(n1399) );
  DFFX1_RVT opC30_d3_reg_4_ ( .D(N1477), .CLK(clk), .QN(n1398) );
  DFFX1_RVT opC30_d3_reg_3_ ( .D(N1476), .CLK(clk), .QN(n1397) );
  DFFX1_RVT opC30_d3_reg_2_ ( .D(N1475), .CLK(clk), .QN(n1396) );
  DFFX1_RVT opC30_d3_reg_1_ ( .D(N1474), .CLK(clk), .QN(n1395) );
  DFFX1_RVT opC30_d3_reg_0_ ( .D(N1473), .CLK(clk), .QN(n1394) );
  DFFX1_RVT opC13_d2_reg_31_ ( .D(N1600), .CLK(clk), .QN(n1297) );
  DFFX1_RVT opC13_d2_reg_30_ ( .D(N1599), .CLK(clk), .QN(n1296) );
  DFFX1_RVT opC13_d2_reg_29_ ( .D(N1598), .CLK(clk), .QN(n1295) );
  DFFX1_RVT opC13_d2_reg_28_ ( .D(N1597), .CLK(clk), .QN(n1294) );
  DFFX1_RVT opC13_d2_reg_27_ ( .D(N1596), .CLK(clk), .QN(n1293) );
  DFFX1_RVT opC13_d2_reg_26_ ( .D(N1595), .CLK(clk), .QN(n1292) );
  DFFX1_RVT opC13_d2_reg_25_ ( .D(N1594), .CLK(clk), .QN(n1291) );
  DFFX1_RVT opC13_d2_reg_24_ ( .D(N1593), .CLK(clk), .QN(n1290) );
  DFFX1_RVT opC13_d2_reg_23_ ( .D(N1592), .CLK(clk), .QN(n1289) );
  DFFX1_RVT opC13_d2_reg_22_ ( .D(N1591), .CLK(clk), .QN(n1288) );
  DFFX1_RVT opC13_d2_reg_21_ ( .D(N1590), .CLK(clk), .QN(n1287) );
  DFFX1_RVT opC13_d2_reg_20_ ( .D(N1589), .CLK(clk), .QN(n1286) );
  DFFX1_RVT opC13_d2_reg_19_ ( .D(N1588), .CLK(clk), .QN(n1285) );
  DFFX1_RVT opC13_d2_reg_18_ ( .D(N1587), .CLK(clk), .QN(n1284) );
  DFFX1_RVT opC13_d2_reg_17_ ( .D(N1586), .CLK(clk), .QN(n1283) );
  DFFX1_RVT opC13_d2_reg_16_ ( .D(N1585), .CLK(clk), .QN(n1282) );
  DFFX1_RVT opC13_d2_reg_15_ ( .D(N1584), .CLK(clk), .QN(n1281) );
  DFFX1_RVT opC13_d2_reg_14_ ( .D(N1583), .CLK(clk), .QN(n1280) );
  DFFX1_RVT opC13_d2_reg_13_ ( .D(N1582), .CLK(clk), .QN(n1279) );
  DFFX1_RVT opC13_d2_reg_12_ ( .D(N1581), .CLK(clk), .QN(n1278) );
  DFFX1_RVT opC13_d2_reg_11_ ( .D(N1580), .CLK(clk), .QN(n1277) );
  DFFX1_RVT opC13_d2_reg_10_ ( .D(N1579), .CLK(clk), .QN(n1276) );
  DFFX1_RVT opC13_d2_reg_9_ ( .D(N1578), .CLK(clk), .QN(n1275) );
  DFFX1_RVT opC13_d2_reg_8_ ( .D(N1577), .CLK(clk), .QN(n1274) );
  DFFX1_RVT opC13_d2_reg_7_ ( .D(N1576), .CLK(clk), .QN(n1273) );
  DFFX1_RVT opC13_d2_reg_6_ ( .D(N1575), .CLK(clk), .QN(n1272) );
  DFFX1_RVT opC13_d2_reg_5_ ( .D(N1574), .CLK(clk), .QN(n1271) );
  DFFX1_RVT opC13_d2_reg_4_ ( .D(N1573), .CLK(clk), .QN(n1270) );
  DFFX1_RVT opC13_d2_reg_3_ ( .D(N1572), .CLK(clk), .QN(n1269) );
  DFFX1_RVT opC13_d2_reg_2_ ( .D(N1571), .CLK(clk), .QN(n1268) );
  DFFX1_RVT opC13_d2_reg_1_ ( .D(N1570), .CLK(clk), .QN(n1267) );
  DFFX1_RVT opC13_d2_reg_0_ ( .D(N1569), .CLK(clk), .QN(n1266) );
  DFFX1_RVT opC22_d2_reg_31_ ( .D(N1664), .CLK(clk), .QN(n1233) );
  DFFX1_RVT opC22_d2_reg_30_ ( .D(N1663), .CLK(clk), .QN(n1232) );
  DFFX1_RVT opC22_d2_reg_29_ ( .D(N1662), .CLK(clk), .QN(n1231) );
  DFFX1_RVT opC22_d2_reg_28_ ( .D(N1661), .CLK(clk), .QN(n1230) );
  DFFX1_RVT opC22_d2_reg_27_ ( .D(N1660), .CLK(clk), .QN(n1229) );
  DFFX1_RVT opC22_d2_reg_26_ ( .D(N1659), .CLK(clk), .QN(n1228) );
  DFFX1_RVT opC22_d2_reg_25_ ( .D(N1658), .CLK(clk), .QN(n1227) );
  DFFX1_RVT opC22_d2_reg_24_ ( .D(N1657), .CLK(clk), .QN(n1226) );
  DFFX1_RVT opC22_d2_reg_23_ ( .D(N1656), .CLK(clk), .QN(n1225) );
  DFFX1_RVT opC22_d2_reg_22_ ( .D(N1655), .CLK(clk), .QN(n1224) );
  DFFX1_RVT opC22_d2_reg_21_ ( .D(N1654), .CLK(clk), .QN(n1223) );
  DFFX1_RVT opC22_d2_reg_20_ ( .D(N1653), .CLK(clk), .QN(n1222) );
  DFFX1_RVT opC22_d2_reg_19_ ( .D(N1652), .CLK(clk), .QN(n1221) );
  DFFX1_RVT opC22_d2_reg_18_ ( .D(N1651), .CLK(clk), .QN(n1220) );
  DFFX1_RVT opC22_d2_reg_17_ ( .D(N1650), .CLK(clk), .QN(n1219) );
  DFFX1_RVT opC22_d2_reg_16_ ( .D(N1649), .CLK(clk), .QN(n1218) );
  DFFX1_RVT opC22_d2_reg_15_ ( .D(N1648), .CLK(clk), .QN(n1217) );
  DFFX1_RVT opC22_d2_reg_14_ ( .D(N1647), .CLK(clk), .QN(n1216) );
  DFFX1_RVT opC22_d2_reg_13_ ( .D(N1646), .CLK(clk), .QN(n1215) );
  DFFX1_RVT opC22_d2_reg_12_ ( .D(N1645), .CLK(clk), .QN(n1214) );
  DFFX1_RVT opC22_d2_reg_11_ ( .D(N1644), .CLK(clk), .QN(n1213) );
  DFFX1_RVT opC22_d2_reg_10_ ( .D(N1643), .CLK(clk), .QN(n1212) );
  DFFX1_RVT opC22_d2_reg_9_ ( .D(N1642), .CLK(clk), .QN(n1211) );
  DFFX1_RVT opC22_d2_reg_8_ ( .D(N1641), .CLK(clk), .QN(n1210) );
  DFFX1_RVT opC22_d2_reg_7_ ( .D(N1640), .CLK(clk), .QN(n1209) );
  DFFX1_RVT opC22_d2_reg_6_ ( .D(N1639), .CLK(clk), .QN(n1208) );
  DFFX1_RVT opC22_d2_reg_5_ ( .D(N1638), .CLK(clk), .QN(n1207) );
  DFFX1_RVT opC22_d2_reg_4_ ( .D(N1637), .CLK(clk), .QN(n1206) );
  DFFX1_RVT opC22_d2_reg_3_ ( .D(N1636), .CLK(clk), .QN(n1205) );
  DFFX1_RVT opC22_d2_reg_2_ ( .D(N1635), .CLK(clk), .QN(n1204) );
  DFFX1_RVT opC22_d2_reg_1_ ( .D(N1634), .CLK(clk), .QN(n1203) );
  DFFX1_RVT opC22_d2_reg_0_ ( .D(N1633), .CLK(clk), .QN(n1202) );
  DFFX1_RVT opC31_d2_reg_31_ ( .D(N1728), .CLK(clk), .QN(n1169) );
  DFFX1_RVT opC31_d2_reg_30_ ( .D(N1727), .CLK(clk), .QN(n1167) );
  DFFX1_RVT opC31_d2_reg_29_ ( .D(N1726), .CLK(clk), .QN(n1165) );
  DFFX1_RVT opC31_d2_reg_28_ ( .D(N1725), .CLK(clk), .QN(n1163) );
  DFFX1_RVT opC31_d2_reg_27_ ( .D(N1724), .CLK(clk), .QN(n1161) );
  DFFX1_RVT opC31_d2_reg_26_ ( .D(N1723), .CLK(clk), .QN(n1159) );
  DFFX1_RVT opC31_d2_reg_25_ ( .D(N1722), .CLK(clk), .QN(n1157) );
  DFFX1_RVT opC31_d2_reg_24_ ( .D(N1721), .CLK(clk), .QN(n1155) );
  DFFX1_RVT opC31_d2_reg_23_ ( .D(N1720), .CLK(clk), .QN(n1153) );
  DFFX1_RVT opC31_d2_reg_22_ ( .D(N1719), .CLK(clk), .QN(n1151) );
  DFFX1_RVT opC31_d2_reg_21_ ( .D(N1718), .CLK(clk), .QN(n1149) );
  DFFX1_RVT opC31_d2_reg_20_ ( .D(N1717), .CLK(clk), .QN(n1147) );
  DFFX1_RVT opC31_d2_reg_19_ ( .D(N1716), .CLK(clk), .QN(n1145) );
  DFFX1_RVT opC31_d2_reg_18_ ( .D(N1715), .CLK(clk), .QN(n1143) );
  DFFX1_RVT opC31_d2_reg_17_ ( .D(N1714), .CLK(clk), .QN(n1141) );
  DFFX1_RVT opC31_d2_reg_16_ ( .D(N1713), .CLK(clk), .QN(n1139) );
  DFFX1_RVT opC31_d2_reg_15_ ( .D(N1712), .CLK(clk), .QN(n1137) );
  DFFX1_RVT opC31_d2_reg_14_ ( .D(N1711), .CLK(clk), .QN(n1135) );
  DFFX1_RVT opC31_d2_reg_13_ ( .D(N1710), .CLK(clk), .QN(n1133) );
  DFFX1_RVT opC31_d2_reg_12_ ( .D(N1709), .CLK(clk), .QN(n1131) );
  DFFX1_RVT opC31_d2_reg_11_ ( .D(N1708), .CLK(clk), .QN(n1129) );
  DFFX1_RVT opC31_d2_reg_10_ ( .D(N1707), .CLK(clk), .QN(n1127) );
  DFFX1_RVT opC31_d2_reg_9_ ( .D(N1706), .CLK(clk), .QN(n1125) );
  DFFX1_RVT opC31_d2_reg_8_ ( .D(N1705), .CLK(clk), .QN(n1123) );
  DFFX1_RVT opC31_d2_reg_7_ ( .D(N1704), .CLK(clk), .QN(n1121) );
  DFFX1_RVT opC31_d2_reg_6_ ( .D(N1703), .CLK(clk), .QN(n1119) );
  DFFX1_RVT opC31_d2_reg_5_ ( .D(N1702), .CLK(clk), .QN(n1117) );
  DFFX1_RVT opC31_d2_reg_4_ ( .D(N1701), .CLK(clk), .QN(n1115) );
  DFFX1_RVT opC31_d2_reg_3_ ( .D(N1700), .CLK(clk), .QN(n1113) );
  DFFX1_RVT opC31_d2_reg_2_ ( .D(N1699), .CLK(clk), .QN(n1111) );
  DFFX1_RVT opC31_d2_reg_1_ ( .D(N1698), .CLK(clk), .QN(n1109) );
  DFFX1_RVT opC31_d2_reg_0_ ( .D(N1697), .CLK(clk), .QN(n1107) );
  DFFX1_RVT opC23_d1_reg_31_ ( .D(N1792), .CLK(clk), .Q(OpC23[31]) );
  DFFX1_RVT opC23_d1_reg_30_ ( .D(N1791), .CLK(clk), .Q(OpC23[30]) );
  DFFX1_RVT opC23_d1_reg_29_ ( .D(N1790), .CLK(clk), .Q(OpC23[29]) );
  DFFX1_RVT opC23_d1_reg_28_ ( .D(N1789), .CLK(clk), .Q(OpC23[28]) );
  DFFX1_RVT opC23_d1_reg_27_ ( .D(N1788), .CLK(clk), .Q(OpC23[27]) );
  DFFX1_RVT opC23_d1_reg_26_ ( .D(N1787), .CLK(clk), .Q(OpC23[26]) );
  DFFX1_RVT opC23_d1_reg_25_ ( .D(N1786), .CLK(clk), .Q(OpC23[25]) );
  DFFX1_RVT opC23_d1_reg_24_ ( .D(N1785), .CLK(clk), .Q(OpC23[24]) );
  DFFX1_RVT opC23_d1_reg_23_ ( .D(N1784), .CLK(clk), .Q(OpC23[23]) );
  DFFX1_RVT opC23_d1_reg_22_ ( .D(N1783), .CLK(clk), .Q(OpC23[22]) );
  DFFX1_RVT opC23_d1_reg_21_ ( .D(N1782), .CLK(clk), .Q(OpC23[21]) );
  DFFX1_RVT opC23_d1_reg_20_ ( .D(N1781), .CLK(clk), .Q(OpC23[20]) );
  DFFX1_RVT opC23_d1_reg_19_ ( .D(N1780), .CLK(clk), .Q(OpC23[19]) );
  DFFX1_RVT opC23_d1_reg_18_ ( .D(N1779), .CLK(clk), .Q(OpC23[18]) );
  DFFX1_RVT opC23_d1_reg_17_ ( .D(N1778), .CLK(clk), .Q(OpC23[17]) );
  DFFX1_RVT opC23_d1_reg_16_ ( .D(N1777), .CLK(clk), .Q(OpC23[16]) );
  DFFX1_RVT opC23_d1_reg_15_ ( .D(N1776), .CLK(clk), .Q(OpC23[15]) );
  DFFX1_RVT opC23_d1_reg_14_ ( .D(N1775), .CLK(clk), .Q(OpC23[14]) );
  DFFX1_RVT opC23_d1_reg_13_ ( .D(N1774), .CLK(clk), .Q(OpC23[13]) );
  DFFX1_RVT opC23_d1_reg_12_ ( .D(N1773), .CLK(clk), .Q(OpC23[12]) );
  DFFX1_RVT opC23_d1_reg_11_ ( .D(N1772), .CLK(clk), .Q(OpC23[11]) );
  DFFX1_RVT opC23_d1_reg_10_ ( .D(N1771), .CLK(clk), .Q(OpC23[10]) );
  DFFX1_RVT opC23_d1_reg_9_ ( .D(N1770), .CLK(clk), .Q(OpC23[9]) );
  DFFX1_RVT opC23_d1_reg_8_ ( .D(N1769), .CLK(clk), .Q(OpC23[8]) );
  DFFX1_RVT opC23_d1_reg_7_ ( .D(N1768), .CLK(clk), .Q(OpC23[7]) );
  DFFX1_RVT opC23_d1_reg_6_ ( .D(N1767), .CLK(clk), .Q(OpC23[6]) );
  DFFX1_RVT opC23_d1_reg_5_ ( .D(N1766), .CLK(clk), .Q(OpC23[5]) );
  DFFX1_RVT opC23_d1_reg_4_ ( .D(N1765), .CLK(clk), .Q(OpC23[4]) );
  DFFX1_RVT opC23_d1_reg_3_ ( .D(N1764), .CLK(clk), .Q(OpC23[3]) );
  DFFX1_RVT opC23_d1_reg_2_ ( .D(N1763), .CLK(clk), .Q(OpC23[2]) );
  DFFX1_RVT opC23_d1_reg_1_ ( .D(N1762), .CLK(clk), .Q(OpC23[1]) );
  DFFX1_RVT opC23_d1_reg_0_ ( .D(N1761), .CLK(clk), .Q(OpC23[0]) );
  DFFX1_RVT opC32_d1_reg_31_ ( .D(N1824), .CLK(clk), .Q(OpC32[31]) );
  DFFX1_RVT opC32_d1_reg_30_ ( .D(N1823), .CLK(clk), .Q(OpC32[30]) );
  DFFX1_RVT opC32_d1_reg_29_ ( .D(N1822), .CLK(clk), .Q(OpC32[29]) );
  DFFX1_RVT opC32_d1_reg_28_ ( .D(N1821), .CLK(clk), .Q(OpC32[28]) );
  DFFX1_RVT opC32_d1_reg_27_ ( .D(N1820), .CLK(clk), .Q(OpC32[27]) );
  DFFX1_RVT opC32_d1_reg_26_ ( .D(N1819), .CLK(clk), .Q(OpC32[26]) );
  DFFX1_RVT opC32_d1_reg_25_ ( .D(N1818), .CLK(clk), .Q(OpC32[25]) );
  DFFX1_RVT opC32_d1_reg_24_ ( .D(N1817), .CLK(clk), .Q(OpC32[24]) );
  DFFX1_RVT opC32_d1_reg_23_ ( .D(N1816), .CLK(clk), .Q(OpC32[23]) );
  DFFX1_RVT opC32_d1_reg_22_ ( .D(N1815), .CLK(clk), .Q(OpC32[22]) );
  DFFX1_RVT opC32_d1_reg_21_ ( .D(N1814), .CLK(clk), .Q(OpC32[21]) );
  DFFX1_RVT opC32_d1_reg_20_ ( .D(N1813), .CLK(clk), .Q(OpC32[20]) );
  DFFX1_RVT opC32_d1_reg_19_ ( .D(N1812), .CLK(clk), .Q(OpC32[19]) );
  DFFX1_RVT opC32_d1_reg_18_ ( .D(N1811), .CLK(clk), .Q(OpC32[18]) );
  DFFX1_RVT opC32_d1_reg_17_ ( .D(N1810), .CLK(clk), .Q(OpC32[17]) );
  DFFX1_RVT opC32_d1_reg_16_ ( .D(N1809), .CLK(clk), .Q(OpC32[16]) );
  DFFX1_RVT opC32_d1_reg_15_ ( .D(N1808), .CLK(clk), .Q(OpC32[15]) );
  DFFX1_RVT opC32_d1_reg_14_ ( .D(N1807), .CLK(clk), .Q(OpC32[14]) );
  DFFX1_RVT opC32_d1_reg_13_ ( .D(N1806), .CLK(clk), .Q(OpC32[13]) );
  DFFX1_RVT opC32_d1_reg_12_ ( .D(N1805), .CLK(clk), .Q(OpC32[12]) );
  DFFX1_RVT opC32_d1_reg_11_ ( .D(N1804), .CLK(clk), .Q(OpC32[11]) );
  DFFX1_RVT opC32_d1_reg_10_ ( .D(N1803), .CLK(clk), .Q(OpC32[10]) );
  DFFX1_RVT opC32_d1_reg_9_ ( .D(N1802), .CLK(clk), .Q(OpC32[9]) );
  DFFX1_RVT opC32_d1_reg_8_ ( .D(N1801), .CLK(clk), .Q(OpC32[8]) );
  DFFX1_RVT opC32_d1_reg_7_ ( .D(N1800), .CLK(clk), .Q(OpC32[7]) );
  DFFX1_RVT opC32_d1_reg_6_ ( .D(N1799), .CLK(clk), .Q(OpC32[6]) );
  DFFX1_RVT opC32_d1_reg_5_ ( .D(N1798), .CLK(clk), .Q(OpC32[5]) );
  DFFX1_RVT opC32_d1_reg_4_ ( .D(N1797), .CLK(clk), .Q(OpC32[4]) );
  DFFX1_RVT opC32_d1_reg_3_ ( .D(N1796), .CLK(clk), .Q(OpC32[3]) );
  DFFX1_RVT opC32_d1_reg_2_ ( .D(N1795), .CLK(clk), .Q(OpC32[2]) );
  DFFX1_RVT opC32_d1_reg_1_ ( .D(N1794), .CLK(clk), .Q(OpC32[1]) );
  DFFX1_RVT opC32_d1_reg_0_ ( .D(N1793), .CLK(clk), .Q(OpC32[0]) );
  DFFSSRX1_RVT opC00_d5_reg_30_ ( .D(1'b0), .SETB(n1075), .RSTB(n3465), .CLK(
        clk), .QN(n3181) );
  DFFSSRX1_RVT opC31_d1_reg_3_ ( .D(1'b0), .SETB(n1113), .RSTB(n3465), .CLK(
        clk), .Q(OpC31[3]) );
  DFFSSRX1_RVT opC11_d4_reg_0_ ( .D(opC11_out[0]), .SETB(1'b1), .RSTB(n3472), 
        .CLK(clk), .QN(n2160) );
  AO22X1_RVT U14 ( .A1(MemOutputB0[66]), .A2(n3540), .A3(MemOutputB0[98]), 
        .A4(n934), .Y(n437) );
  AO22X1_RVT U16 ( .A1(MemOutputB0[68]), .A2(n3540), .A3(MemOutputB0[100]), 
        .A4(n935), .Y(n421) );
  AOI22X1_RVT U49 ( .A1(MemOutputB0[211]), .A2(n3504), .A3(MemOutputB0[243]), 
        .A4(n3331), .Y(n403) );
  AO22X1_RVT U189 ( .A1(n3533), .A2(MemOutputB0[77]), .A3(MemOutputB0[109]), 
        .A4(n3236), .Y(n509) );
  AO22X1_RVT U253 ( .A1(MemOutputA0[68]), .A2(n3542), .A3(MemOutputA0[100]), 
        .A4(n3236), .Y(n933) );
  AO22X1_RVT U274 ( .A1(MemOutputB0[74]), .A2(n3241), .A3(MemOutputB0[106]), 
        .A4(n3236), .Y(n521) );
  AO22X1_RVT U344 ( .A1(MemOutputA0[74]), .A2(n3541), .A3(MemOutputA0[106]), 
        .A4(n3521), .Y(n1033) );
  AO22X1_RVT U478 ( .A1(MemOutputA3[71]), .A2(n3541), .A3(MemOutputA3[103]), 
        .A4(n3508), .Y(n537) );
  NBUFFX2_RVT U494 ( .A(n3290), .Y(n3291) );
  AO22X2_RVT U530 ( .A1(MemOutputB0[78]), .A2(n3540), .A3(MemOutputB0[110]), 
        .A4(n3236), .Y(n505) );
  AO22X2_RVT U531 ( .A1(MemOutputB0[79]), .A2(n3540), .A3(MemOutputB0[111]), 
        .A4(n3515), .Y(n501) );
  AO22X2_RVT U533 ( .A1(MemOutputB0[94]), .A2(n3542), .A3(MemOutputB0[126]), 
        .A4(n3523), .Y(n433) );
  AO22X2_RVT U534 ( .A1(MemOutputA3[70]), .A2(n3539), .A3(MemOutputA3[102]), 
        .A4(n3523), .Y(n541) );
  AO22X2_RVT U535 ( .A1(MemOutputB0[71]), .A2(n3542), .A3(MemOutputB0[103]), 
        .A4(n3523), .Y(n409) );
  DELLN3X2_RVT U536 ( .A(n934), .Y(n3517) );
  DELLN3X2_RVT U538 ( .A(n934), .Y(n3507) );
  DELLN3X2_RVT U539 ( .A(n934), .Y(n3512) );
  DELLN3X2_RVT U540 ( .A(n935), .Y(n3506) );
  DELLN3X2_RVT U541 ( .A(n935), .Y(n3519) );
  DELLN3X2_RVT U542 ( .A(n935), .Y(n3510) );
  AO22X2_RVT U543 ( .A1(MemOutputB0[95]), .A2(n3541), .A3(MemOutputB0[127]), 
        .A4(n3522), .Y(n429) );
  DELLN3X2_RVT U544 ( .A(n3522), .Y(n3518) );
  DELLN3X2_RVT U545 ( .A(n3522), .Y(n3509) );
  DELLN2X2_RVT U555 ( .A(n3522), .Y(n3520) );
  DELLN3X2_RVT U556 ( .A(n3522), .Y(n3511) );
  DELLN1X2_RVT U557 ( .A(n1034), .Y(n12) );
  NAND3X0_RVT U558 ( .A1(n1), .A2(n4), .A3(n5), .Y(ipA0[5]) );
  AOI22X1_RVT U559 ( .A1(MemOutputA0[197]), .A2(n3501), .A3(MemOutputA0[229]), 
        .A4(n3322), .Y(n1) );
  AOI22X1_RVT U567 ( .A1(MemOutputA0[165]), .A2(n3248), .A3(MemOutputA0[133]), 
        .A4(n3272), .Y(n4) );
  AOI221X1_RVT U570 ( .A1(MemOutputA0[5]), .A2(n3291), .A3(MemOutputA0[37]), 
        .A4(n3561), .A5(n929), .Y(n5) );
  IBUFFX2_RVT U572 ( .A(n3565), .Y(n3293) );
  NBUFFX2_RVT U574 ( .A(n471), .Y(n3282) );
  IBUFFX2_RVT U575 ( .A(n484), .Y(n10) );
  IBUFFX2_RVT U577 ( .A(n9), .Y(n3565) );
  IBUFFX2_RVT U580 ( .A(n484), .Y(n3562) );
  DELLN1X2_RVT U581 ( .A(n455), .Y(n3324) );
  DELLN3X2_RVT U583 ( .A(n3335), .Y(n3330) );
  DELLN3X2_RVT U584 ( .A(n3335), .Y(n3332) );
  DELLN3X2_RVT U585 ( .A(n3335), .Y(n3334) );
  DELLN2X2_RVT U586 ( .A(n3335), .Y(n3327) );
  DELLN3X2_RVT U588 ( .A(n3309), .Y(n3319) );
  INVX0_RVT U589 ( .A(latCnt[1]), .Y(n936) );
  IBUFFX2_RVT U590 ( .A(n3242), .Y(n3268) );
  IBUFFX2_RVT U591 ( .A(n3540), .Y(n14) );
  IBUFFX4_RVT U593 ( .A(n14), .Y(n15) );
  NBUFFX2_RVT U594 ( .A(n3273), .Y(n3278) );
  AOI22X1_RVT U595 ( .A1(MemOutputB0[201]), .A2(n3492), .A3(MemOutputB0[233]), 
        .A4(n3310), .Y(n407) );
  AOI22X1_RVT U596 ( .A1(MemOutputB0[171]), .A2(n3254), .A3(MemOutputB0[139]), 
        .A4(n3287), .Y(n474) );
  NBUFFX2_RVT U598 ( .A(n3302), .Y(n3304) );
  NBUFFX2_RVT U599 ( .A(n471), .Y(n3270) );
  NBUFFX2_RVT U600 ( .A(n456), .Y(n3303) );
  AO22X1_RVT U601 ( .A1(MemOutputA3[203]), .A2(n3495), .A3(MemOutputA3[235]), 
        .A4(n3318), .Y(n642) );
  INVX0_RVT U603 ( .A(n3566), .Y(n3292) );
  NBUFFX2_RVT U604 ( .A(n3292), .Y(n3305) );
  NBUFFX2_RVT U605 ( .A(n3269), .Y(n3271) );
  NBUFFX2_RVT U606 ( .A(n3268), .Y(n3288) );
  INVX0_RVT U608 ( .A(n3569), .Y(n3482) );
  NBUFFX2_RVT U609 ( .A(n3287), .Y(n3283) );
  IBUFFX2_RVT U610 ( .A(n3566), .Y(n456) );
  IBUFFX2_RVT U611 ( .A(n3483), .Y(n3309) );
  DELLN1X2_RVT U613 ( .A(n3269), .Y(n3273) );
  NBUFFX2_RVT U614 ( .A(n3301), .Y(n3298) );
  DELLN2X2_RVT U615 ( .A(n3269), .Y(n3272) );
  DELLN1X2_RVT U616 ( .A(n506), .Y(n454) );
  NAND3X0_RVT U618 ( .A1(n16), .A2(n398), .A3(n399), .Y(ipB0[8]) );
  AOI22X1_RVT U619 ( .A1(MemOutputB0[200]), .A2(n3492), .A3(MemOutputB0[232]), 
        .A4(n3329), .Y(n16) );
  AOI22X1_RVT U620 ( .A1(MemOutputB0[168]), .A2(n3266), .A3(MemOutputB0[136]), 
        .A4(n3270), .Y(n398) );
  AOI221X1_RVT U621 ( .A1(MemOutputB0[8]), .A2(n3301), .A3(MemOutputB0[40]), 
        .A4(n10), .A5(n405), .Y(n399) );
  DELLN1X2_RVT U623 ( .A(n3299), .Y(n3296) );
  INVX0_RVT U624 ( .A(latCnt[2]), .Y(n3571) );
  IBUFFX2_RVT U625 ( .A(n3242), .Y(n470) );
  INVX0_RVT U626 ( .A(latCnt[0]), .Y(n947) );
  INVX0_RVT U628 ( .A(latCnt[3]), .Y(n486) );
  INVX0_RVT U629 ( .A(n491), .Y(n3503) );
  NAND3X0_RVT U635 ( .A1(n3237), .A2(n3238), .A3(n3239), .Y(ipB0[27]) );
  AO22X1_RVT U636 ( .A1(MemOutputA3[194]), .A2(n3493), .A3(MemOutputA3[226]), 
        .A4(n3319), .Y(n562) );
  AO22X1_RVT U638 ( .A1(MemOutputB1[208]), .A2(n3491), .A3(MemOutputB1[240]), 
        .A4(n3320), .Y(n366) );
  NBUFFX2_RVT U639 ( .A(n3547), .Y(n3551) );
  NBUFFX2_RVT U640 ( .A(n3271), .Y(n3281) );
  NBUFFX2_RVT U641 ( .A(n3317), .Y(n3313) );
  NBUFFX2_RVT U643 ( .A(n3316), .Y(n3312) );
  NBUFFX2_RVT U644 ( .A(n3278), .Y(n3276) );
  AO22X1_RVT U645 ( .A1(MemOutputA3[190]), .A2(n3248), .A3(MemOutputA3[158]), 
        .A4(n3288), .Y(n559) );
  AO22X1_RVT U646 ( .A1(MemOutputB2[206]), .A2(n3488), .A3(MemOutputB2[238]), 
        .A4(n3320), .Y(n246) );
  AO22X1_RVT U648 ( .A1(MemOutputB2[219]), .A2(n3487), .A3(MemOutputB2[251]), 
        .A4(n3319), .Y(n190) );
  AO22X1_RVT U649 ( .A1(MemOutputA1[192]), .A2(n3500), .A3(MemOutputA1[224]), 
        .A4(n3319), .Y(n906) );
  AO22X1_RVT U650 ( .A1(MemOutputA1[169]), .A2(n3249), .A3(MemOutputA1[137]), 
        .A4(n454), .Y(n783) );
  IBUFFX2_RVT U651 ( .A(n3240), .Y(n3244) );
  NBUFFX2_RVT U653 ( .A(n17), .Y(n455) );
  INVX0_RVT U654 ( .A(n3267), .Y(n3544) );
  INVX0_RVT U655 ( .A(n3267), .Y(n3543) );
  OR3X2_RVT U656 ( .A1(n434), .A2(n435), .A3(n436), .Y(ipB0[2]) );
  NBUFFX2_RVT U657 ( .A(n3276), .Y(n506) );
  NBUFFX2_RVT U658 ( .A(n3243), .Y(n3249) );
  INVX0_RVT U659 ( .A(n17), .Y(n3483) );
  NBUFFX2_RVT U660 ( .A(n3330), .Y(n3317) );
  OR3X2_RVT U661 ( .A1(n1022), .A2(n1023), .A3(n1024), .Y(ipA0[12]) );
  OR3X2_RVT U662 ( .A1(n1014), .A2(n1015), .A3(n1016), .Y(ipA0[14]) );
  OR3X2_RVT U663 ( .A1(n1018), .A2(n1019), .A3(n1020), .Y(ipA0[13]) );
  NBUFFX2_RVT U664 ( .A(n3564), .Y(n3547) );
  IBUFFX2_RVT U665 ( .A(n450), .Y(n451) );
  NBUFFX2_RVT U666 ( .A(n514), .Y(n3262) );
  OR3X2_RVT U667 ( .A1(n918), .A2(n919), .A3(n920), .Y(ipA0[7]) );
  NBUFFX2_RVT U668 ( .A(n3506), .Y(n3508) );
  NBUFFX2_RVT U669 ( .A(n3332), .Y(n3316) );
  INVX0_RVT U670 ( .A(n3267), .Y(n507) );
  INVX0_RVT U671 ( .A(n3267), .Y(n519) );
  OR3X1_RVT U673 ( .A1(n430), .A2(n431), .A3(n432), .Y(ipB0[30]) );
  NAND3X0_RVT U674 ( .A1(n400), .A2(n402), .A3(n403), .Y(ipB0[19]) );
  AOI221X1_RVT U675 ( .A1(MemOutputB0[19]), .A2(n3293), .A3(MemOutputB0[51]), 
        .A4(n10), .A5(n485), .Y(n400) );
  AOI22X1_RVT U676 ( .A1(MemOutputB0[179]), .A2(n3266), .A3(MemOutputB0[147]), 
        .A4(n452), .Y(n402) );
  AOI22X1_RVT U678 ( .A1(MemOutputB0[203]), .A2(n3504), .A3(MemOutputB0[235]), 
        .A4(n3311), .Y(n472) );
  NBUFFX2_RVT U679 ( .A(n456), .Y(n3308) );
  NAND3X0_RVT U680 ( .A1(n404), .A2(n406), .A3(n407), .Y(ipB0[9]) );
  AOI221X1_RVT U681 ( .A1(MemOutputB0[9]), .A2(n456), .A3(MemOutputB0[41]), 
        .A4(n3564), .A5(n401), .Y(n404) );
  AOI22X1_RVT U682 ( .A1(MemOutputB0[169]), .A2(n3253), .A3(MemOutputB0[137]), 
        .A4(n3279), .Y(n406) );
  NBUFFX2_RVT U683 ( .A(n3290), .Y(n408) );
  DELLN3X2_RVT U684 ( .A(n3309), .Y(n3320) );
  NBUFFX2_RVT U685 ( .A(n456), .Y(n3307) );
  OR3X2_RVT U686 ( .A1(n914), .A2(n915), .A3(n916), .Y(ipA0[8]) );
  NAND3X0_RVT U688 ( .A1(n418), .A2(n419), .A3(n420), .Y(ipB0[10]) );
  AOI22X1_RVT U689 ( .A1(MemOutputB0[202]), .A2(n3492), .A3(MemOutputB0[234]), 
        .A4(n3326), .Y(n418) );
  AOI22X1_RVT U702 ( .A1(MemOutputB0[170]), .A2(n3261), .A3(MemOutputB0[138]), 
        .A4(n3275), .Y(n419) );
  AOI221X1_RVT U707 ( .A1(MemOutputB0[10]), .A2(n456), .A3(MemOutputB0[42]), 
        .A4(n3553), .A5(n521), .Y(n420) );
  NBUFFX2_RVT U733 ( .A(n3542), .Y(n3539) );
  NAND3X0_RVT U739 ( .A1(n438), .A2(n439), .A3(n440), .Y(ipB0[4]) );
  AOI22X1_RVT U839 ( .A1(MemOutputB0[196]), .A2(n3492), .A3(MemOutputB0[228]), 
        .A4(n3310), .Y(n438) );
  AOI22X1_RVT U948 ( .A1(MemOutputB0[164]), .A2(n3251), .A3(MemOutputB0[132]), 
        .A4(n3285), .Y(n439) );
  AOI221X1_RVT U1009 ( .A1(MemOutputB0[4]), .A2(n456), .A3(MemOutputB0[36]), 
        .A4(n10), .A5(n421), .Y(n440) );
  NAND3X0_RVT U1013 ( .A1(n442), .A2(n443), .A3(n444), .Y(ipB0[7]) );
  AOI22X1_RVT U1073 ( .A1(MemOutputB0[199]), .A2(n3492), .A3(MemOutputB0[231]), 
        .A4(n3322), .Y(n442) );
  AOI22X1_RVT U1169 ( .A1(MemOutputB0[167]), .A2(n3252), .A3(MemOutputB0[135]), 
        .A4(n3282), .Y(n443) );
  AOI221X1_RVT U1175 ( .A1(MemOutputB0[7]), .A2(n3302), .A3(MemOutputB0[39]), 
        .A4(n3562), .A5(n409), .Y(n444) );
  OR3X2_RVT U1180 ( .A1(n922), .A2(n923), .A3(n924), .Y(ipA0[6]) );
  AO22X1_RVT U1185 ( .A1(MemOutputB1[179]), .A2(n3258), .A3(MemOutputB1[147]), 
        .A4(n3282), .Y(n355) );
  AO22X1_RVT U1190 ( .A1(MemOutputB2[190]), .A2(n3252), .A3(MemOutputB2[158]), 
        .A4(n3283), .Y(n175) );
  AO22X1_RVT U1191 ( .A1(MemOutputA0[176]), .A2(n3252), .A3(MemOutputA0[144]), 
        .A4(n3277), .Y(n1007) );
  IBUFFX2_RVT U1193 ( .A(n3240), .Y(n3255) );
  INVX0_RVT U1194 ( .A(latCnt[1]), .Y(n3570) );
  NBUFFX2_RVT U1195 ( .A(n1034), .Y(n3540) );
  OR3X2_RVT U1196 ( .A1(n1030), .A2(n1031), .A3(n1032), .Y(ipA0[10]) );
  AND4X1_RVT U1197 ( .A1(latCnt[0]), .A2(n3572), .A3(latCnt[1]), .A4(latCnt[2]), .Y(n17) );
  NBUFFX2_RVT U1198 ( .A(n1034), .Y(n3241) );
  AO22X2_RVT U1199 ( .A1(MemOutputA2[180]), .A2(n3253), .A3(MemOutputA2[148]), 
        .A4(n3277), .Y(n731) );
  AO22X2_RVT U1200 ( .A1(MemOutputA1[187]), .A2(n3263), .A3(MemOutputA1[155]), 
        .A4(n3282), .Y(n831) );
  AND4X1_RVT U1215 ( .A1(n947), .A2(n936), .A3(n3571), .A4(n948), .Y(n9) );
  INVX0_RVT U1216 ( .A(latCnt[3]), .Y(n948) );
  IBUFFX2_RVT U1218 ( .A(n3256), .Y(n450) );
  NBUFFX2_RVT U1219 ( .A(n470), .Y(n452) );
  INVX0_RVT U1270 ( .A(n3565), .Y(n3294) );
  NBUFFX2_RVT U1271 ( .A(n500), .Y(n3246) );
  NBUFFX2_RVT U1272 ( .A(n3290), .Y(n3306) );
  IBUFFX2_RVT U1273 ( .A(n9), .Y(n3566) );
  NAND3X0_RVT U1274 ( .A1(n458), .A2(n459), .A3(n460), .Y(ipB0[17]) );
  AOI221X1_RVT U1293 ( .A1(MemOutputB0[17]), .A2(n3301), .A3(MemOutputB0[49]), 
        .A4(n3562), .A5(n493), .Y(n458) );
  AOI22X1_RVT U1300 ( .A1(MemOutputB0[177]), .A2(n3256), .A3(MemOutputB0[145]), 
        .A4(n3274), .Y(n459) );
  AOI22X2_RVT U1305 ( .A1(MemOutputB0[209]), .A2(n3502), .A3(MemOutputB0[241]), 
        .A4(n3311), .Y(n460) );
  NBUFFX2_RVT U1310 ( .A(n514), .Y(n3263) );
  OR3X1_RVT U1320 ( .A1(n412), .A2(n411), .A3(n410), .Y(ipB0[6]) );
  NBUFFX2_RVT U1322 ( .A(n3300), .Y(n3295) );
  NBUFFX2_RVT U1325 ( .A(n3295), .Y(n3297) );
  NBUFFX2_RVT U1326 ( .A(n3540), .Y(n3541) );
  AOI22X1_RVT U1328 ( .A1(MemOutputB0[205]), .A2(n3502), .A3(MemOutputB0[237]), 
        .A4(n3321), .Y(n466) );
  NAND3X0_RVT U1329 ( .A1(n462), .A2(n463), .A3(n464), .Y(ipB0[24]) );
  AOI221X1_RVT U1330 ( .A1(n3306), .A2(MemOutputB0[24]), .A3(MemOutputB0[56]), 
        .A4(n3564), .A5(n461), .Y(n462) );
  AOI22X1_RVT U1331 ( .A1(MemOutputB0[184]), .A2(n3243), .A3(MemOutputB0[152]), 
        .A4(n3280), .Y(n463) );
  AOI22X1_RVT U1332 ( .A1(MemOutputB0[216]), .A2(n3504), .A3(MemOutputB0[248]), 
        .A4(n3321), .Y(n464) );
  NAND3X0_RVT U1333 ( .A1(n466), .A2(n467), .A3(n468), .Y(ipB0[13]) );
  AOI22X1_RVT U1334 ( .A1(MemOutputB0[173]), .A2(n3244), .A3(MemOutputB0[141]), 
        .A4(n3274), .Y(n467) );
  AOI221X1_RVT U1335 ( .A1(MemOutputB0[13]), .A2(n3292), .A3(MemOutputB0[45]), 
        .A4(n3553), .A5(n509), .Y(n468) );
  IBUFFX2_RVT U1336 ( .A(n3242), .Y(n471) );
  NAND3X0_RVT U1337 ( .A1(n472), .A2(n474), .A3(n475), .Y(ipB0[11]) );
  AOI221X1_RVT U1338 ( .A1(MemOutputB0[11]), .A2(n3293), .A3(MemOutputB0[43]), 
        .A4(n3553), .A5(n517), .Y(n475) );
  NAND3X0_RVT U1339 ( .A1(n476), .A2(n482), .A3(n483), .Y(ipB0[12]) );
  AOI22X1_RVT U1340 ( .A1(MemOutputB0[204]), .A2(n3502), .A3(MemOutputB0[236]), 
        .A4(n3331), .Y(n476) );
  AOI22X2_RVT U1341 ( .A1(MemOutputB0[172]), .A2(n3246), .A3(MemOutputB0[140]), 
        .A4(n3287), .Y(n482) );
  AOI221X1_RVT U1374 ( .A1(MemOutputB0[12]), .A2(n3292), .A3(MemOutputB0[44]), 
        .A4(n3553), .A5(n513), .Y(n483) );
  NAND4X1_RVT U1794 ( .A1(n520), .A2(n3570), .A3(n3571), .A4(n486), .Y(n484)
         );
  AO22X2_RVT U2844 ( .A1(MemOutputB3[205]), .A2(n3486), .A3(MemOutputB3[237]), 
        .A4(n3309), .Y(n122) );
  AO22X2_RVT U2846 ( .A1(MemOutputA2[192]), .A2(n3497), .A3(MemOutputA2[224]), 
        .A4(n3309), .Y(n778) );
  AOI22X2_RVT U2847 ( .A1(MemOutputB0[219]), .A2(n3502), .A3(MemOutputB0[251]), 
        .A4(n3309), .Y(n3237) );
  NAND3X0_RVT U2848 ( .A1(n502), .A2(n503), .A3(n504), .Y(ipB0[15]) );
  NAND3X0_RVT U2849 ( .A1(n487), .A2(n488), .A3(n490), .Y(ipA0[3]) );
  AOI22X2_RVT U2850 ( .A1(MemOutputA0[195]), .A2(n3501), .A3(MemOutputA0[227]), 
        .A4(n3333), .Y(n487) );
  AOI221X1_RVT U2851 ( .A1(MemOutputA0[3]), .A2(n408), .A3(MemOutputA0[35]), 
        .A4(n10), .A5(n937), .Y(n488) );
  AOI22X1_RVT U2852 ( .A1(MemOutputA0[163]), .A2(n3266), .A3(MemOutputA0[131]), 
        .A4(n3287), .Y(n490) );
  NAND4X1_RVT U2853 ( .A1(n948), .A2(n947), .A3(latCnt[1]), .A4(latCnt[2]), 
        .Y(n491) );
  NAND3X0_RVT U2854 ( .A1(n492), .A2(n494), .A3(n495), .Y(ipA0[4]) );
  AOI221X1_RVT U2855 ( .A1(MemOutputA0[4]), .A2(n456), .A3(MemOutputA0[36]), 
        .A4(n3562), .A5(n933), .Y(n492) );
  AOI22X1_RVT U2856 ( .A1(MemOutputA0[164]), .A2(n3251), .A3(MemOutputA0[132]), 
        .A4(n3279), .Y(n494) );
  AOI22X1_RVT U2857 ( .A1(MemOutputA0[196]), .A2(n3501), .A3(MemOutputA0[228]), 
        .A4(n3324), .Y(n495) );
  NAND3X0_RVT U2858 ( .A1(n496), .A2(n498), .A3(n499), .Y(ipB0[14]) );
  AOI221X1_RVT U2859 ( .A1(MemOutputB0[14]), .A2(n3301), .A3(MemOutputB0[46]), 
        .A4(n3553), .A5(n505), .Y(n496) );
  AOI22X1_RVT U2860 ( .A1(MemOutputB0[174]), .A2(n3244), .A3(MemOutputB0[142]), 
        .A4(n452), .Y(n498) );
  AOI22X1_RVT U2861 ( .A1(MemOutputB0[206]), .A2(n3505), .A3(MemOutputB0[238]), 
        .A4(n3309), .Y(n499) );
  IBUFFX2_RVT U2862 ( .A(n3240), .Y(n500) );
  NBUFFX2_RVT U2863 ( .A(n3261), .Y(n514) );
  NAND3X0_RVT U2864 ( .A1(n930), .A2(n931), .A3(n932), .Y(ipB0[26]) );
  INVX0_RVT U2865 ( .A(latCnt[3]), .Y(n3572) );
  AOI22X1_RVT U2866 ( .A1(MemOutputB0[207]), .A2(n3505), .A3(MemOutputB0[239]), 
        .A4(n3309), .Y(n502) );
  AOI22X1_RVT U2867 ( .A1(MemOutputB0[175]), .A2(n3246), .A3(MemOutputB0[143]), 
        .A4(n3274), .Y(n503) );
  AOI221X1_RVT U2868 ( .A1(MemOutputB0[15]), .A2(n408), .A3(MemOutputB0[47]), 
        .A4(n3553), .A5(n501), .Y(n504) );
  NBUFFX2_RVT U2869 ( .A(n17), .Y(n3335) );
  INVX0_RVT U2870 ( .A(n3566), .Y(n3300) );
  NBUFFX2_RVT U2871 ( .A(n13), .Y(n508) );
  NAND3X0_RVT U2872 ( .A1(n512), .A2(n511), .A3(n510), .Y(ipB0[25]) );
  AOI221X1_RVT U2873 ( .A1(MemOutputB0[25]), .A2(n408), .A3(MemOutputB0[57]), 
        .A4(n3562), .A5(n457), .Y(n510) );
  AOI22X1_RVT U2874 ( .A1(MemOutputB0[185]), .A2(n3244), .A3(MemOutputB0[153]), 
        .A4(n3284), .Y(n511) );
  AOI22X1_RVT U2875 ( .A1(MemOutputB0[217]), .A2(n3504), .A3(MemOutputB0[249]), 
        .A4(n3328), .Y(n512) );
  NAND3X0_RVT U2876 ( .A1(n515), .A2(n516), .A3(n518), .Y(ipB0[22]) );
  AOI22X1_RVT U2877 ( .A1(MemOutputB0[214]), .A2(n3504), .A3(MemOutputB0[246]), 
        .A4(n3331), .Y(n515) );
  AOI22X1_RVT U2878 ( .A1(MemOutputB0[182]), .A2(n3245), .A3(MemOutputB0[150]), 
        .A4(n3269), .Y(n516) );
  AOI221X1_RVT U2879 ( .A1(MemOutputB0[22]), .A2(n3294), .A3(MemOutputB0[54]), 
        .A4(n3564), .A5(n469), .Y(n518) );
  IBUFFX2_RVT U2880 ( .A(n3539), .Y(n3267) );
  NBUFFX2_RVT U2881 ( .A(latCnt[0]), .Y(n520) );
  NAND3X0_RVT U2882 ( .A1(n522), .A2(n523), .A3(n524), .Y(ipB0[21]) );
  AOI22X1_RVT U2883 ( .A1(MemOutputB0[213]), .A2(n3505), .A3(MemOutputB0[245]), 
        .A4(n3331), .Y(n522) );
  AOI22X1_RVT U2884 ( .A1(MemOutputB0[181]), .A2(n3243), .A3(MemOutputB0[149]), 
        .A4(n3284), .Y(n523) );
  AOI221X1_RVT U2885 ( .A1(MemOutputB0[21]), .A2(n3300), .A3(MemOutputB0[53]), 
        .A4(n10), .A5(n473), .Y(n524) );
  NAND3X0_RVT U2886 ( .A1(n928), .A2(n927), .A3(n926), .Y(ipB0[20]) );
  AOI221X1_RVT U2887 ( .A1(MemOutputB0[20]), .A2(n3300), .A3(MemOutputB0[52]), 
        .A4(n10), .A5(n477), .Y(n926) );
  AOI22X1_RVT U2888 ( .A1(MemOutputB0[180]), .A2(n3243), .A3(MemOutputB0[148]), 
        .A4(n471), .Y(n927) );
  AOI22X1_RVT U2889 ( .A1(MemOutputB0[212]), .A2(n3502), .A3(MemOutputB0[244]), 
        .A4(n3331), .Y(n928) );
  DELLN2X2_RVT U2890 ( .A(n3562), .Y(n3548) );
  DELLN2X2_RVT U2891 ( .A(n3564), .Y(n3549) );
  DELLN2X2_RVT U2892 ( .A(n3562), .Y(n3550) );
  INVX0_RVT U2893 ( .A(latCnt[2]), .Y(n946) );
  NBUFFX2_RVT U2894 ( .A(n13), .Y(n3514) );
  AOI221X1_RVT U2895 ( .A1(MemOutputB0[26]), .A2(n3293), .A3(MemOutputB0[58]), 
        .A4(n3562), .A5(n453), .Y(n930) );
  AOI22X1_RVT U2896 ( .A1(MemOutputB0[186]), .A2(n3266), .A3(MemOutputB0[154]), 
        .A4(n452), .Y(n931) );
  AOI22X1_RVT U2897 ( .A1(MemOutputB0[218]), .A2(n3502), .A3(MemOutputB0[250]), 
        .A4(n3321), .Y(n932) );
  AND4X1_RVT U2898 ( .A1(n948), .A2(n946), .A3(n947), .A4(latCnt[1]), .Y(n1034) );
  IBUFFX2_RVT U2899 ( .A(n3524), .Y(n934) );
  IBUFFX2_RVT U2900 ( .A(n3524), .Y(n935) );
  IBUFFX2_RVT U2901 ( .A(n3524), .Y(n3522) );
  NBUFFX2_RVT U2902 ( .A(n13), .Y(n3515) );
  NAND3X0_RVT U2903 ( .A1(n3227), .A2(n3228), .A3(n3229), .Y(ipA0[2]) );
  IBUFFX2_RVT U2904 ( .A(n3524), .Y(n3523) );
  IBUFFX2_RVT U2905 ( .A(n491), .Y(n3502) );
  IBUFFX2_RVT U2906 ( .A(n491), .Y(n3505) );
  IBUFFX2_RVT U2907 ( .A(n491), .Y(n3504) );
  AOI22X1_RVT U2908 ( .A1(MemOutputB0[188]), .A2(n3260), .A3(MemOutputB0[156]), 
        .A4(n3286), .Y(n991) );
  NAND3X0_RVT U2909 ( .A1(n990), .A2(n991), .A3(n992), .Y(ipB0[28]) );
  AOI22X1_RVT U2910 ( .A1(MemOutputB0[220]), .A2(n3492), .A3(MemOutputB0[252]), 
        .A4(n3336), .Y(n990) );
  AOI221X1_RVT U2911 ( .A1(MemOutputB0[28]), .A2(n408), .A3(MemOutputB0[60]), 
        .A4(n10), .A5(n445), .Y(n992) );
  IBUFFX2_RVT U2912 ( .A(n484), .Y(n3563) );
  IBUFFX2_RVT U2913 ( .A(n484), .Y(n3564) );
  IBUFFX2_RVT U2914 ( .A(n13), .Y(n3524) );
  OR3X2_RVT U2915 ( .A1(n1035), .A2(n1036), .A3(n1038), .Y(ipB0[0]) );
  AO22X1_RVT U2916 ( .A1(MemOutputB0[192]), .A2(n3484), .A3(MemOutputB0[224]), 
        .A4(n3334), .Y(n1035) );
  AO22X1_RVT U2917 ( .A1(MemOutputB0[160]), .A2(n3264), .A3(MemOutputB0[128]), 
        .A4(n452), .Y(n1036) );
  AO221X1_RVT U2918 ( .A1(MemOutputB0[0]), .A2(n408), .A3(MemOutputB0[32]), 
        .A4(n3552), .A5(n525), .Y(n1038) );
  NBUFFX2_RVT U2919 ( .A(n3464), .Y(n3373) );
  NBUFFX2_RVT U2920 ( .A(n3464), .Y(n3374) );
  NBUFFX2_RVT U2921 ( .A(n3464), .Y(n3375) );
  NBUFFX2_RVT U2922 ( .A(n3463), .Y(n3376) );
  NBUFFX2_RVT U2923 ( .A(n3463), .Y(n3377) );
  NBUFFX2_RVT U2924 ( .A(n3463), .Y(n3378) );
  NBUFFX2_RVT U2925 ( .A(n3462), .Y(n3379) );
  NBUFFX2_RVT U2926 ( .A(n3462), .Y(n3380) );
  NBUFFX2_RVT U2927 ( .A(n3461), .Y(n3382) );
  NBUFFX2_RVT U2928 ( .A(n3461), .Y(n3383) );
  NBUFFX2_RVT U2929 ( .A(n3461), .Y(n3384) );
  NBUFFX2_RVT U2930 ( .A(n3460), .Y(n3385) );
  NBUFFX2_RVT U2931 ( .A(n3460), .Y(n3386) );
  NBUFFX2_RVT U2932 ( .A(n3460), .Y(n3387) );
  NBUFFX2_RVT U2933 ( .A(n3459), .Y(n3388) );
  NBUFFX2_RVT U2934 ( .A(n3459), .Y(n3389) );
  NBUFFX2_RVT U2935 ( .A(n3459), .Y(n3390) );
  NBUFFX2_RVT U2936 ( .A(n3458), .Y(n3391) );
  NBUFFX2_RVT U2937 ( .A(n3458), .Y(n3392) );
  NBUFFX2_RVT U2938 ( .A(n3457), .Y(n3393) );
  NBUFFX2_RVT U2939 ( .A(n3457), .Y(n3395) );
  NBUFFX2_RVT U2940 ( .A(n3456), .Y(n3396) );
  NBUFFX2_RVT U2941 ( .A(n3456), .Y(n3397) );
  NBUFFX2_RVT U2942 ( .A(n3456), .Y(n3398) );
  NBUFFX2_RVT U2943 ( .A(n3455), .Y(n3399) );
  NBUFFX2_RVT U2944 ( .A(n3455), .Y(n3400) );
  NBUFFX2_RVT U2945 ( .A(n3455), .Y(n3401) );
  NBUFFX2_RVT U2946 ( .A(n3454), .Y(n3402) );
  NBUFFX2_RVT U2947 ( .A(n3454), .Y(n3403) );
  NBUFFX2_RVT U2948 ( .A(n3454), .Y(n3404) );
  NBUFFX2_RVT U2949 ( .A(n3453), .Y(n3405) );
  NBUFFX2_RVT U2950 ( .A(n3453), .Y(n3406) );
  NBUFFX2_RVT U2951 ( .A(n3453), .Y(n3407) );
  NBUFFX2_RVT U2952 ( .A(n3457), .Y(n3394) );
  NBUFFX2_RVT U2953 ( .A(n3463), .Y(n3408) );
  NBUFFX2_RVT U2954 ( .A(n3461), .Y(n3409) );
  NBUFFX2_RVT U2955 ( .A(n3462), .Y(n3410) );
  NBUFFX2_RVT U2956 ( .A(n3459), .Y(n3411) );
  NBUFFX2_RVT U2957 ( .A(n3458), .Y(n3412) );
  NBUFFX2_RVT U2958 ( .A(n3459), .Y(n3413) );
  NBUFFX2_RVT U2959 ( .A(n3452), .Y(n3414) );
  NBUFFX2_RVT U2960 ( .A(n3452), .Y(n3415) );
  NBUFFX2_RVT U2961 ( .A(n3452), .Y(n3416) );
  NBUFFX2_RVT U2962 ( .A(n3451), .Y(n3417) );
  NBUFFX2_RVT U2963 ( .A(n3462), .Y(n3381) );
  NBUFFX2_RVT U2964 ( .A(n3451), .Y(n3419) );
  NBUFFX2_RVT U2965 ( .A(n3450), .Y(n3420) );
  NBUFFX2_RVT U2966 ( .A(n3450), .Y(n3421) );
  NBUFFX2_RVT U2967 ( .A(n3449), .Y(n3423) );
  NBUFFX2_RVT U2968 ( .A(n3449), .Y(n3424) );
  NBUFFX2_RVT U2969 ( .A(n3449), .Y(n3425) );
  NBUFFX2_RVT U2970 ( .A(n3448), .Y(n3426) );
  NBUFFX2_RVT U2971 ( .A(n3450), .Y(n3422) );
  NBUFFX2_RVT U2972 ( .A(n3448), .Y(n3427) );
  NBUFFX2_RVT U2973 ( .A(n3448), .Y(n3428) );
  NBUFFX2_RVT U2974 ( .A(n3447), .Y(n3429) );
  NBUFFX2_RVT U2975 ( .A(n3447), .Y(n3430) );
  NBUFFX2_RVT U2976 ( .A(n3447), .Y(n3431) );
  NBUFFX2_RVT U2977 ( .A(n3446), .Y(n3432) );
  NBUFFX2_RVT U2978 ( .A(n3446), .Y(n3433) );
  NBUFFX2_RVT U2979 ( .A(n3446), .Y(n3434) );
  NBUFFX2_RVT U2980 ( .A(n3445), .Y(n3435) );
  NBUFFX2_RVT U2981 ( .A(n3451), .Y(n3418) );
  NBUFFX2_RVT U2982 ( .A(n3445), .Y(n3436) );
  NBUFFX2_RVT U2983 ( .A(n3444), .Y(n3437) );
  NBUFFX2_RVT U2984 ( .A(n3444), .Y(n3438) );
  NBUFFX2_RVT U2985 ( .A(n3443), .Y(n3439) );
  NBUFFX2_RVT U2986 ( .A(n3443), .Y(n3440) );
  NBUFFX2_RVT U2987 ( .A(n3465), .Y(n3372) );
  NBUFFX2_RVT U2988 ( .A(n3468), .Y(n3362) );
  NBUFFX2_RVT U2989 ( .A(n3468), .Y(n3361) );
  NBUFFX2_RVT U2990 ( .A(n3468), .Y(n3360) );
  NBUFFX2_RVT U2991 ( .A(n3468), .Y(n3363) );
  NBUFFX2_RVT U2992 ( .A(n3467), .Y(n3366) );
  NBUFFX2_RVT U2993 ( .A(n3467), .Y(n3365) );
  NBUFFX2_RVT U2994 ( .A(n3467), .Y(n3364) );
  NBUFFX2_RVT U2995 ( .A(n3473), .Y(n3367) );
  NBUFFX2_RVT U2996 ( .A(n3479), .Y(n3370) );
  NBUFFX2_RVT U2997 ( .A(n3467), .Y(n3369) );
  NBUFFX2_RVT U2998 ( .A(n3478), .Y(n3368) );
  NBUFFX2_RVT U2999 ( .A(n3470), .Y(n3371) );
  NBUFFX2_RVT U3000 ( .A(n3468), .Y(n3359) );
  NBUFFX2_RVT U3001 ( .A(n3468), .Y(n3343) );
  NBUFFX2_RVT U3002 ( .A(n3480), .Y(n3347) );
  NBUFFX2_RVT U3003 ( .A(n3481), .Y(n3346) );
  NBUFFX2_RVT U3004 ( .A(n3471), .Y(n3345) );
  NBUFFX2_RVT U3005 ( .A(n3471), .Y(n3351) );
  NBUFFX2_RVT U3006 ( .A(n3471), .Y(n3350) );
  NBUFFX2_RVT U3007 ( .A(n3469), .Y(n3344) );
  NBUFFX2_RVT U3008 ( .A(n3471), .Y(n3349) );
  NBUFFX2_RVT U3009 ( .A(n3478), .Y(n3348) );
  NBUFFX2_RVT U3010 ( .A(n3468), .Y(n3358) );
  NBUFFX2_RVT U3011 ( .A(n3470), .Y(n3353) );
  NBUFFX2_RVT U3012 ( .A(n3470), .Y(n3352) );
  NBUFFX2_RVT U3013 ( .A(n3469), .Y(n3357) );
  NBUFFX2_RVT U3014 ( .A(n3469), .Y(n3356) );
  NBUFFX2_RVT U3015 ( .A(n3469), .Y(n3355) );
  NBUFFX2_RVT U3016 ( .A(n3470), .Y(n3354) );
  NBUFFX2_RVT U3017 ( .A(n3442), .Y(n3441) );
  NBUFFX2_RVT U3018 ( .A(n3482), .Y(n3468) );
  NBUFFX2_RVT U3019 ( .A(n3473), .Y(n3467) );
  NBUFFX2_RVT U3020 ( .A(n3473), .Y(n3466) );
  NBUFFX2_RVT U3021 ( .A(n3473), .Y(n3471) );
  NBUFFX2_RVT U3022 ( .A(n3473), .Y(n3469) );
  NBUFFX2_RVT U3023 ( .A(n3473), .Y(n3470) );
  NBUFFX2_RVT U3024 ( .A(n3482), .Y(n3465) );
  NBUFFX2_RVT U3025 ( .A(n3482), .Y(n3464) );
  NBUFFX2_RVT U3026 ( .A(n3474), .Y(n3463) );
  NBUFFX2_RVT U3027 ( .A(n3474), .Y(n3461) );
  NBUFFX2_RVT U3028 ( .A(n3475), .Y(n3460) );
  NBUFFX2_RVT U3029 ( .A(n3475), .Y(n3459) );
  NBUFFX2_RVT U3030 ( .A(n3475), .Y(n3458) );
  NBUFFX2_RVT U3031 ( .A(n3476), .Y(n3456) );
  NBUFFX2_RVT U3032 ( .A(n3476), .Y(n3455) );
  NBUFFX2_RVT U3033 ( .A(n3477), .Y(n3454) );
  NBUFFX2_RVT U3034 ( .A(n3477), .Y(n3453) );
  NBUFFX2_RVT U3035 ( .A(n3476), .Y(n3457) );
  NBUFFX2_RVT U3036 ( .A(n3478), .Y(n3452) );
  NBUFFX2_RVT U3037 ( .A(n3474), .Y(n3462) );
  NBUFFX2_RVT U3038 ( .A(n3479), .Y(n3449) );
  NBUFFX2_RVT U3039 ( .A(n3479), .Y(n3450) );
  NBUFFX2_RVT U3040 ( .A(n3479), .Y(n3448) );
  NBUFFX2_RVT U3041 ( .A(n3480), .Y(n3447) );
  NBUFFX2_RVT U3042 ( .A(n3480), .Y(n3446) );
  NBUFFX2_RVT U3043 ( .A(n3478), .Y(n3451) );
  NBUFFX2_RVT U3044 ( .A(n3481), .Y(n3444) );
  NBUFFX2_RVT U3045 ( .A(n3481), .Y(n3443) );
  NBUFFX2_RVT U3046 ( .A(n3481), .Y(n3442) );
  NBUFFX2_RVT U3047 ( .A(n3480), .Y(n3445) );
  NBUFFX2_RVT U3048 ( .A(n3477), .Y(n3472) );
  NBUFFX2_RVT U3049 ( .A(n507), .Y(n3525) );
  NBUFFX2_RVT U3050 ( .A(n519), .Y(n3526) );
  NBUFFX2_RVT U3051 ( .A(n3544), .Y(n3530) );
  NBUFFX2_RVT U3052 ( .A(n3544), .Y(n3529) );
  NBUFFX2_RVT U3053 ( .A(n3544), .Y(n3531) );
  NBUFFX2_RVT U3054 ( .A(n3543), .Y(n3537) );
  NBUFFX2_RVT U3055 ( .A(n3543), .Y(n3536) );
  NBUFFX2_RVT U3056 ( .A(n3543), .Y(n3538) );
  NBUFFX2_RVT U3057 ( .A(n3554), .Y(n3560) );
  NBUFFX2_RVT U3058 ( .A(n3544), .Y(n3527) );
  NBUFFX2_RVT U3059 ( .A(n3544), .Y(n3528) );
  NBUFFX2_RVT U3060 ( .A(n3543), .Y(n3534) );
  NBUFFX2_RVT U3061 ( .A(n3543), .Y(n3535) );
  NBUFFX2_RVT U3062 ( .A(n3482), .Y(n3473) );
  NBUFFX2_RVT U3063 ( .A(rstnPipe), .Y(n3475) );
  NBUFFX2_RVT U3064 ( .A(n3482), .Y(n3476) );
  NBUFFX2_RVT U3065 ( .A(n3482), .Y(n3477) );
  NBUFFX2_RVT U3066 ( .A(rstnPipe), .Y(n3474) );
  NBUFFX2_RVT U3067 ( .A(n3482), .Y(n3479) );
  NBUFFX2_RVT U3068 ( .A(n3482), .Y(n3478) );
  NBUFFX2_RVT U3069 ( .A(n3482), .Y(n3481) );
  NBUFFX2_RVT U3070 ( .A(n3482), .Y(n3480) );
  NBUFFX2_RVT U3071 ( .A(n3563), .Y(n3553) );
  NBUFFX2_RVT U3072 ( .A(n3562), .Y(n3545) );
  NBUFFX2_RVT U3073 ( .A(n3564), .Y(n3546) );
  NBUFFX2_RVT U3074 ( .A(n3563), .Y(n3552) );
  NBUFFX2_RVT U3075 ( .A(n3506), .Y(n3516) );
  NBUFFX2_RVT U3076 ( .A(n3507), .Y(n3513) );
  NBUFFX2_RVT U3077 ( .A(n3502), .Y(n3497) );
  NBUFFX2_RVT U3078 ( .A(n3503), .Y(n3501) );
  NBUFFX2_RVT U3079 ( .A(n3505), .Y(n3500) );
  NBUFFX2_RVT U3080 ( .A(n3560), .Y(n3559) );
  NBUFFX2_RVT U3081 ( .A(n3550), .Y(n3557) );
  NBUFFX2_RVT U3082 ( .A(n3560), .Y(n3558) );
  NBUFFX2_RVT U3083 ( .A(n3504), .Y(n3488) );
  NBUFFX2_RVT U3084 ( .A(n3504), .Y(n3490) );
  NBUFFX2_RVT U3085 ( .A(n3504), .Y(n3489) );
  NBUFFX2_RVT U3086 ( .A(n3550), .Y(n3555) );
  NBUFFX2_RVT U3087 ( .A(n3554), .Y(n3556) );
  NBUFFX2_RVT U3088 ( .A(n3499), .Y(n3491) );
  NBUFFX2_RVT U3089 ( .A(n3502), .Y(n3494) );
  NBUFFX2_RVT U3090 ( .A(n3502), .Y(n3495) );
  NBUFFX2_RVT U3091 ( .A(n3485), .Y(n3499) );
  NBUFFX2_RVT U3092 ( .A(n3504), .Y(n3486) );
  NBUFFX2_RVT U3093 ( .A(n3504), .Y(n3487) );
  NBUFFX2_RVT U3094 ( .A(n3505), .Y(n3485) );
  NBUFFX2_RVT U3095 ( .A(n3505), .Y(n3484) );
  NBUFFX2_RVT U3096 ( .A(n3499), .Y(n3493) );
  NBUFFX2_RVT U3097 ( .A(n3514), .Y(n3521) );
  NBUFFX2_RVT U3098 ( .A(n1034), .Y(n3532) );
  NBUFFX2_RVT U3099 ( .A(n1034), .Y(n3533) );
  INVX1_RVT U3100 ( .A(rstnPipe), .Y(n3567) );
  INVX1_RVT U3101 ( .A(rstnPipe), .Y(n3568) );
  INVX1_RVT U3102 ( .A(n3), .Y(n3573) );
  INVX1_RVT U3103 ( .A(rstnPipe), .Y(n3569) );
  INVX1_RVT U3104 ( .A(addrInc), .Y(n3574) );
  NAND3X0_RVT U3105 ( .A1(n1039), .A2(n1040), .A3(n1041), .Y(ipB0[16]) );
  AOI22X1_RVT U3106 ( .A1(MemOutputB0[208]), .A2(n3505), .A3(MemOutputB0[240]), 
        .A4(n3311), .Y(n1039) );
  AOI22X1_RVT U3107 ( .A1(MemOutputB0[176]), .A2(n3246), .A3(MemOutputB0[144]), 
        .A4(n3274), .Y(n1040) );
  AOI221X1_RVT U3108 ( .A1(MemOutputB0[16]), .A2(n3293), .A3(MemOutputB0[48]), 
        .A4(n3553), .A5(n497), .Y(n1041) );
  NAND3X0_RVT U3109 ( .A1(n1112), .A2(n3180), .A3(n3226), .Y(ipB0[23]) );
  AOI22X1_RVT U3110 ( .A1(MemOutputB0[215]), .A2(n3504), .A3(MemOutputB0[247]), 
        .A4(n3328), .Y(n1112) );
  AOI22X1_RVT U3111 ( .A1(MemOutputB0[183]), .A2(n3244), .A3(MemOutputB0[151]), 
        .A4(n3268), .Y(n3180) );
  AOI221X1_RVT U3112 ( .A1(MemOutputB0[23]), .A2(n3293), .A3(MemOutputB0[55]), 
        .A4(n10), .A5(n465), .Y(n3226) );
  AOI22X1_RVT U3113 ( .A1(MemOutputA0[194]), .A2(n3502), .A3(MemOutputA0[226]), 
        .A4(n3321), .Y(n3227) );
  AOI22X1_RVT U3114 ( .A1(MemOutputA0[162]), .A2(n3256), .A3(MemOutputA0[130]), 
        .A4(n3284), .Y(n3228) );
  AOI221X1_RVT U3115 ( .A1(MemOutputA0[2]), .A2(n3300), .A3(MemOutputA0[34]), 
        .A4(n3562), .A5(n949), .Y(n3229) );
  AO22X1_RVT U3116 ( .A1(MemOutputB0[222]), .A2(n3492), .A3(MemOutputB0[254]), 
        .A4(n3324), .Y(n430) );
  NAND3X0_RVT U3117 ( .A1(n3230), .A2(n3231), .A3(n3232), .Y(ipB0[18]) );
  AOI22X1_RVT U3118 ( .A1(MemOutputB0[210]), .A2(n3505), .A3(MemOutputB0[242]), 
        .A4(n3311), .Y(n3230) );
  AOI22X1_RVT U3119 ( .A1(MemOutputB0[178]), .A2(n3244), .A3(MemOutputB0[146]), 
        .A4(n3284), .Y(n3231) );
  AOI221X1_RVT U3120 ( .A1(MemOutputB0[18]), .A2(n3292), .A3(MemOutputB0[50]), 
        .A4(n10), .A5(n489), .Y(n3232) );
  NAND3X0_RVT U3121 ( .A1(n3233), .A2(n3234), .A3(n3235), .Y(ipA0[1]) );
  AOI22X1_RVT U3122 ( .A1(MemOutputA0[193]), .A2(n3505), .A3(MemOutputA0[225]), 
        .A4(n3328), .Y(n3233) );
  AOI22X1_RVT U3123 ( .A1(MemOutputA0[161]), .A2(n3244), .A3(MemOutputA0[129]), 
        .A4(n3280), .Y(n3234) );
  AOI221X1_RVT U3124 ( .A1(n3306), .A2(MemOutputA0[1]), .A3(MemOutputA0[33]), 
        .A4(n3564), .A5(n993), .Y(n3235) );
  AOI22X1_RVT U3125 ( .A1(MemOutputB0[221]), .A2(n3492), .A3(MemOutputB0[253]), 
        .A4(n3325), .Y(n3340) );
  AND4X1_RVT U3126 ( .A1(n486), .A2(n946), .A3(n520), .A4(latCnt[1]), .Y(n13)
         );
  NAND3X0_RVT U3127 ( .A1(n3337), .A2(n3338), .A3(n3339), .Y(ipA0[0]) );
  AO22X1_RVT U3128 ( .A1(n12), .A2(MemOutputA0[65]), .A3(n3514), .A4(
        MemOutputA0[97]), .Y(n993) );
  NBUFFX2_RVT U3129 ( .A(n3502), .Y(n3498) );
  NBUFFX2_RVT U3130 ( .A(n3502), .Y(n3496) );
  NAND3X0_RVT U3131 ( .A1(n3340), .A2(n3341), .A3(n3342), .Y(ipB0[29]) );
  IBUFFX2_RVT U3132 ( .A(n3240), .Y(n3245) );
  IBUFFX2_RVT U3133 ( .A(n3240), .Y(n3243) );
  IBUFFX2_RVT U3134 ( .A(n3242), .Y(n3269) );
  NBUFFX2_RVT U3135 ( .A(n1034), .Y(n3542) );
  NBUFFX2_RVT U3136 ( .A(n3548), .Y(n3554) );
  NBUFFX2_RVT U3137 ( .A(n3563), .Y(n3561) );
  NBUFFX2_RVT U3138 ( .A(n13), .Y(n3236) );
  AOI22X1_RVT U3139 ( .A1(MemOutputB0[187]), .A2(n3243), .A3(MemOutputB0[155]), 
        .A4(n3280), .Y(n3238) );
  AOI221X1_RVT U3140 ( .A1(MemOutputB0[27]), .A2(n3291), .A3(MemOutputB0[59]), 
        .A4(n10), .A5(n449), .Y(n3239) );
  NAND4X1_RVT U3141 ( .A1(n486), .A2(n936), .A3(n520), .A4(latCnt[2]), .Y(
        n3240) );
  NAND4X1_RVT U3142 ( .A1(n486), .A2(n3570), .A3(n947), .A4(latCnt[2]), .Y(
        n3242) );
  NBUFFX2_RVT U3143 ( .A(n3503), .Y(n3492) );
  NBUFFX2_RVT U3144 ( .A(n3245), .Y(n3247) );
  NBUFFX2_RVT U3145 ( .A(n3245), .Y(n3248) );
  NBUFFX2_RVT U3146 ( .A(n500), .Y(n3250) );
  NBUFFX2_RVT U3147 ( .A(n3244), .Y(n3251) );
  NBUFFX2_RVT U3148 ( .A(n500), .Y(n3252) );
  NBUFFX2_RVT U3149 ( .A(n3244), .Y(n3253) );
  NBUFFX2_RVT U3150 ( .A(n500), .Y(n3254) );
  NBUFFX2_RVT U3151 ( .A(n3255), .Y(n3256) );
  NBUFFX2_RVT U3152 ( .A(n3243), .Y(n3257) );
  NBUFFX2_RVT U3153 ( .A(n500), .Y(n3258) );
  NBUFFX2_RVT U3154 ( .A(n3243), .Y(n3259) );
  NBUFFX2_RVT U3155 ( .A(n3245), .Y(n3260) );
  NBUFFX2_RVT U3156 ( .A(n3255), .Y(n3261) );
  NBUFFX2_RVT U3157 ( .A(n3243), .Y(n3264) );
  NBUFFX2_RVT U3158 ( .A(n3247), .Y(n3265) );
  NBUFFX2_RVT U3159 ( .A(n3245), .Y(n3266) );
  NBUFFX2_RVT U3160 ( .A(n3269), .Y(n3274) );
  NBUFFX2_RVT U3161 ( .A(n3268), .Y(n3275) );
  NBUFFX2_RVT U3162 ( .A(n3269), .Y(n3277) );
  NBUFFX2_RVT U3163 ( .A(n3268), .Y(n3279) );
  NBUFFX2_RVT U3164 ( .A(n470), .Y(n3280) );
  NBUFFX2_RVT U3165 ( .A(n470), .Y(n3284) );
  NBUFFX2_RVT U3166 ( .A(n3268), .Y(n3285) );
  NBUFFX2_RVT U3167 ( .A(n471), .Y(n3286) );
  NBUFFX2_RVT U3168 ( .A(n471), .Y(n3287) );
  NBUFFX2_RVT U3169 ( .A(n508), .Y(n3289) );
  NBUFFX2_RVT U3170 ( .A(n9), .Y(n3290) );
  NBUFFX2_RVT U3171 ( .A(n456), .Y(n3299) );
  NBUFFX2_RVT U3172 ( .A(n3290), .Y(n3301) );
  NBUFFX2_RVT U3173 ( .A(n3294), .Y(n3302) );
  NBUFFX2_RVT U3174 ( .A(n3335), .Y(n3310) );
  NBUFFX2_RVT U3175 ( .A(n455), .Y(n3311) );
  NBUFFX2_RVT U3176 ( .A(n3311), .Y(n3314) );
  NBUFFX2_RVT U3177 ( .A(n3309), .Y(n3315) );
  NBUFFX2_RVT U3178 ( .A(n3309), .Y(n3318) );
  NBUFFX2_RVT U3179 ( .A(n455), .Y(n3321) );
  NBUFFX2_RVT U3180 ( .A(n3335), .Y(n3322) );
  NBUFFX2_RVT U3181 ( .A(n3335), .Y(n3323) );
  NBUFFX2_RVT U3182 ( .A(n3335), .Y(n3325) );
  NBUFFX2_RVT U3183 ( .A(n455), .Y(n3326) );
  NBUFFX2_RVT U3184 ( .A(n455), .Y(n3328) );
  NBUFFX2_RVT U3185 ( .A(n3335), .Y(n3329) );
  NBUFFX2_RVT U3186 ( .A(n455), .Y(n3331) );
  NBUFFX2_RVT U3187 ( .A(n455), .Y(n3333) );
  NBUFFX2_RVT U3188 ( .A(n3335), .Y(n3336) );
  AOI22X1_RVT U3189 ( .A1(MemOutputA0[192]), .A2(n3505), .A3(MemOutputA0[224]), 
        .A4(n3328), .Y(n3337) );
  AOI22X1_RVT U3190 ( .A1(MemOutputA0[160]), .A2(n3243), .A3(MemOutputA0[128]), 
        .A4(n3280), .Y(n3338) );
  AOI221X1_RVT U3191 ( .A1(MemOutputA0[0]), .A2(n3306), .A3(MemOutputA0[32]), 
        .A4(n3562), .A5(n1037), .Y(n3339) );
  AOI22X1_RVT U3192 ( .A1(MemOutputB0[189]), .A2(n3246), .A3(MemOutputB0[157]), 
        .A4(n3287), .Y(n3341) );
  AOI221X1_RVT U3193 ( .A1(MemOutputB0[29]), .A2(n3292), .A3(MemOutputB0[61]), 
        .A4(n10), .A5(n441), .Y(n3342) );
endmodule


module TOP ( clk, rstnSys, startSys, MemOutputA0, MemOutputA1, MemOutputA2, 
        MemOutputA3, MemOutputB0, MemOutputB1, MemOutputB2, MemOutputB3, OpC00, 
        OpC01, OpC02, OpC03, OpC10, OpC11, OpC12, OpC13, OpC20, OpC21, OpC22, 
        OpC23, OpC30, OpC31, OpC32, OpC33, BankAddr, start_check );
  input [255:0] MemOutputA0;
  input [255:0] MemOutputA1;
  input [255:0] MemOutputA2;
  input [255:0] MemOutputA3;
  input [255:0] MemOutputB0;
  input [255:0] MemOutputB1;
  input [255:0] MemOutputB2;
  input [255:0] MemOutputB3;
  output [31:0] OpC00;
  output [31:0] OpC01;
  output [31:0] OpC02;
  output [31:0] OpC03;
  output [31:0] OpC10;
  output [31:0] OpC11;
  output [31:0] OpC12;
  output [31:0] OpC13;
  output [31:0] OpC20;
  output [31:0] OpC21;
  output [31:0] OpC22;
  output [31:0] OpC23;
  output [31:0] OpC30;
  output [31:0] OpC31;
  output [31:0] OpC32;
  output [31:0] OpC33;
  output [9:0] BankAddr;
  input clk, rstnSys, startSys;
  output start_check;
  wire   rstnPipe, rstnAddr, addrInc;
  wire   [15:0] rstnPsum;
  wire   [3:0] latCnt;

  CTRL ctrl ( .clk(clk), .rstnSys(rstnSys), .startSys(startSys), .rstnPsum(
        rstnPsum), .rstnPipe(rstnPipe), .rstnAddr(rstnAddr), .addrInc(addrInc), 
        .latCnt(latCnt), .start_check(start_check) );
  DATA data ( .clk(clk), .rstnPipe(rstnPipe), .rstnAddr(rstnAddr), .addrInc(
        addrInc), .rstnPsum(rstnPsum), .latCnt(latCnt), .MemOutputA0(
        MemOutputA0), .MemOutputA1(MemOutputA1), .MemOutputA2(MemOutputA2), 
        .MemOutputA3(MemOutputA3), .MemOutputB0(MemOutputB0), .MemOutputB1(
        MemOutputB1), .MemOutputB2(MemOutputB2), .MemOutputB3(MemOutputB3), 
        .OpC00(OpC00), .OpC01(OpC01), .OpC02(OpC02), .OpC03(OpC03), .OpC10(
        OpC10), .OpC11(OpC11), .OpC12(OpC12), .OpC13(OpC13), .OpC20(OpC20), 
        .OpC21(OpC21), .OpC22(OpC22), .OpC23(OpC23), .OpC30(OpC30), .OpC31(
        OpC31), .OpC32(OpC32), .OpC33(OpC33), .BankAddr(BankAddr) );
endmodule

